-------------------------------------------------------------------------------
-- Title      : Slow ADC Look-up-tables for the environmental data conversion
-- Project    : EPIX Detector
-------------------------------------------------------------------------------
-- File       : SlowAdcLUT.vhd
-- Company    : SLAC National Accelerator Laboratory
-------------------------------------------------------------------------------
-- Description:
-- This block is responsible for the conversion of the voltages, currents
-- temperatures from the ADS1217 to the human readable data
-------------------------------------------------------------------------------
-- This file is part of 'EPIX Development Firmware'.
-- It is subject to the license terms in the LICENSE.txt file found in the
-- top-level directory of this distribution and at:
--    https://confluence.slac.stanford.edu/display/ppareg/LICENSE.html.
-- No part of 'EPIX Development Firmware', including this file,
-- may be copied, modified, propagated, or distributed except according to
-- the terms contained in the LICENSE.txt file.
-------------------------------------------------------------------------------

LIBRARY ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library surf;
use surf.StdRtlPkg.all;

library epix_hr_core;
use epix_hr_core.SlowAdcPkg.all;

--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--
library unisim;
use unisim.vcomponents.all;

entity SlowAdcLUT is
   port (
      -- Master system clock
      sysClk          : in  std_logic;
      sysClkRst       : in  std_logic;

      -- ADC raw data inputs
      adcData         : in Slv24Array(8 downto 0);

      -- Converted data outputs
      outEnvData      : out Slv32Array(8 downto 0)
   );
end SlowAdcLUT;


-- Define architecture
architecture RTL of SlowAdcLUT is

   signal th0_address_a :     std_logic_vector(15 downto 0);
   signal th0_h_data_out_a :  std_logic_vector(35 downto 0);
   signal th0_l_data_out_a :  std_logic_vector(35 downto 0);
   signal th0_data_out_a :    std_logic_vector(15 downto 0);

   signal th1_address_a :     std_logic_vector(15 downto 0);
   signal th1_h_data_out_a :  std_logic_vector(35 downto 0);
   signal th1_l_data_out_a :  std_logic_vector(35 downto 0);
   signal th1_data_out_a :    std_logic_vector(15 downto 0);

   signal hum_address_a :     std_logic_vector(15 downto 0);
   signal hum_h_data_out_a :  std_logic_vector(35 downto 0);
   signal hum_l_data_out_a :  std_logic_vector(35 downto 0);
   signal hum_data_out_a :    std_logic_vector(15 downto 0);

   signal iana_address_a :    std_logic_vector(15 downto 0);
   signal iana_h_data_out_a : std_logic_vector(35 downto 0);
   signal iana_l_data_out_a : std_logic_vector(35 downto 0);

   signal idig_address_a :    std_logic_vector(15 downto 0);
   signal idig_h_data_out_a : std_logic_vector(35 downto 0);
   signal idig_l_data_out_a : std_logic_vector(35 downto 0);

   signal igua_address_a :    std_logic_vector(15 downto 0);
   signal igua_h_data_out_a : std_logic_vector(35 downto 0);
   signal igua_l_data_out_a : std_logic_vector(35 downto 0);

   signal ibia_address_a :    std_logic_vector(15 downto 0);
   signal ibia_h_data_out_a : std_logic_vector(35 downto 0);
   signal ibia_l_data_out_a : std_logic_vector(35 downto 0);

   signal avin_address_a :    std_logic_vector(15 downto 0);
   signal avin_h_data_out_a : std_logic_vector(35 downto 0);
   signal avin_l_data_out_a : std_logic_vector(35 downto 0);

   signal dvin_address_a :    std_logic_vector(15 downto 0);
   signal dvin_h_data_out_a : std_logic_vector(35 downto 0);
   signal dvin_l_data_out_a : std_logic_vector(35 downto 0);

begin


   th0_h_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_H_TH0_00,
      INIT_01 => INIT_H_TH0_01,
      INIT_02 => INIT_H_TH0_02,
      INIT_03 => INIT_H_TH0_03,
      INIT_04 => INIT_H_TH0_04,
      INIT_05 => INIT_H_TH0_05,
      INIT_06 => INIT_H_TH0_06,
      INIT_07 => INIT_H_TH0_07,
      INIT_08 => INIT_H_TH0_08,
      INIT_09 => INIT_H_TH0_09,
      INIT_0A => INIT_H_TH0_0A,
      INIT_0B => INIT_H_TH0_0B,
      INIT_0C => INIT_H_TH0_0C,
      INIT_0D => INIT_H_TH0_0D,
      INIT_0E => INIT_H_TH0_0E,
      INIT_0F => INIT_H_TH0_0F,
      INIT_10 => INIT_H_TH0_10,
      INIT_11 => INIT_H_TH0_11,
      INIT_12 => INIT_H_TH0_12,
      INIT_13 => INIT_H_TH0_13,
      INIT_14 => INIT_H_TH0_14,
      INIT_15 => INIT_H_TH0_15,
      INIT_16 => INIT_H_TH0_16,
      INIT_17 => INIT_H_TH0_17,
      INIT_18 => INIT_H_TH0_18,
      INIT_19 => INIT_H_TH0_19,
      INIT_1A => INIT_H_TH0_1A,
      INIT_1B => INIT_H_TH0_1B,
      INIT_1C => INIT_H_TH0_1C,
      INIT_1D => INIT_H_TH0_1D,
      INIT_1E => INIT_H_TH0_1E,
      INIT_1F => INIT_H_TH0_1F,
      INIT_20 => INIT_H_TH0_20,
      INIT_21 => INIT_H_TH0_21,
      INIT_22 => INIT_H_TH0_22,
      INIT_23 => INIT_H_TH0_23,
      INIT_24 => INIT_H_TH0_24,
      INIT_25 => INIT_H_TH0_25,
      INIT_26 => INIT_H_TH0_26,
      INIT_27 => INIT_H_TH0_27,
      INIT_28 => INIT_H_TH0_28,
      INIT_29 => INIT_H_TH0_29,
      INIT_2A => INIT_H_TH0_2A,
      INIT_2B => INIT_H_TH0_2B,
      INIT_2C => INIT_H_TH0_2C,
      INIT_2D => INIT_H_TH0_2D,
      INIT_2E => INIT_H_TH0_2E,
      INIT_2F => INIT_H_TH0_2F,
      INIT_30 => INIT_H_TH0_30,
      INIT_31 => INIT_H_TH0_31,
      INIT_32 => INIT_H_TH0_32,
      INIT_33 => INIT_H_TH0_33,
      INIT_34 => INIT_H_TH0_34,
      INIT_35 => INIT_H_TH0_35,
      INIT_36 => INIT_H_TH0_36,
      INIT_37 => INIT_H_TH0_37,
      INIT_38 => INIT_H_TH0_38,
      INIT_39 => INIT_H_TH0_39,
      INIT_3A => INIT_H_TH0_3A,
      INIT_3B => INIT_H_TH0_3B,
      INIT_3C => INIT_H_TH0_3C,
      INIT_3D => INIT_H_TH0_3D,
      INIT_3E => INIT_H_TH0_3E,
      INIT_3F => INIT_H_TH0_3F,
      INIT_40 => INIT_H_TH0_40,
      INIT_41 => INIT_H_TH0_41,
      INIT_42 => INIT_H_TH0_42,
      INIT_43 => INIT_H_TH0_43,
      INIT_44 => INIT_H_TH0_44,
      INIT_45 => INIT_H_TH0_45,
      INIT_46 => INIT_H_TH0_46,
      INIT_47 => INIT_H_TH0_47,
      INIT_48 => INIT_H_TH0_48,
      INIT_49 => INIT_H_TH0_49,
      INIT_4A => INIT_H_TH0_4A,
      INIT_4B => INIT_H_TH0_4B,
      INIT_4C => INIT_H_TH0_4C,
      INIT_4D => INIT_H_TH0_4D,
      INIT_4E => INIT_H_TH0_4E,
      INIT_4F => INIT_H_TH0_4F,
      INIT_50 => INIT_H_TH0_50,
      INIT_51 => INIT_H_TH0_51,
      INIT_52 => INIT_H_TH0_52,
      INIT_53 => INIT_H_TH0_53,
      INIT_54 => INIT_H_TH0_54,
      INIT_55 => INIT_H_TH0_55,
      INIT_56 => INIT_H_TH0_56,
      INIT_57 => INIT_H_TH0_57,
      INIT_58 => INIT_H_TH0_58,
      INIT_59 => INIT_H_TH0_59,
      INIT_5A => INIT_H_TH0_5A,
      INIT_5B => INIT_H_TH0_5B,
      INIT_5C => INIT_H_TH0_5C,
      INIT_5D => INIT_H_TH0_5D,
      INIT_5E => INIT_H_TH0_5E,
      INIT_5F => INIT_H_TH0_5F,
      INIT_60 => INIT_H_TH0_60,
      INIT_61 => INIT_H_TH0_61,
      INIT_62 => INIT_H_TH0_62,
      INIT_63 => INIT_H_TH0_63,
      INIT_64 => INIT_H_TH0_64,
      INIT_65 => INIT_H_TH0_65,
      INIT_66 => INIT_H_TH0_66,
      INIT_67 => INIT_H_TH0_67,
      INIT_68 => INIT_H_TH0_68,
      INIT_69 => INIT_H_TH0_69,
      INIT_6A => INIT_H_TH0_6A,
      INIT_6B => INIT_H_TH0_6B,
      INIT_6C => INIT_H_TH0_6C,
      INIT_6D => INIT_H_TH0_6D,
      INIT_6E => INIT_H_TH0_6E,
      INIT_6F => INIT_H_TH0_6F,
      INIT_70 => INIT_H_TH0_70,
      INIT_71 => INIT_H_TH0_71,
      INIT_72 => INIT_H_TH0_72,
      INIT_73 => INIT_H_TH0_73,
      INIT_74 => INIT_H_TH0_74,
      INIT_75 => INIT_H_TH0_75,
      INIT_76 => INIT_H_TH0_76,
      INIT_77 => INIT_H_TH0_77,
      INIT_78 => INIT_H_TH0_78,
      INIT_79 => INIT_H_TH0_79,
      INIT_7A => INIT_H_TH0_7A,
      INIT_7B => INIT_H_TH0_7B,
      INIT_7C => INIT_H_TH0_7C,
      INIT_7D => INIT_H_TH0_7D,
      INIT_7E => INIT_H_TH0_7E,
      INIT_7F => INIT_H_TH0_7F
   ) port map(
      ADDRARDADDR    => th0_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => th0_h_data_out_a(31 downto 0),
      DOPADOP        => th0_h_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );



   th0_l_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_L_TH0_00,
      INIT_01 => INIT_L_TH0_01,
      INIT_02 => INIT_L_TH0_02,
      INIT_03 => INIT_L_TH0_03,
      INIT_04 => INIT_L_TH0_04,
      INIT_05 => INIT_L_TH0_05,
      INIT_06 => INIT_L_TH0_06,
      INIT_07 => INIT_L_TH0_07,
      INIT_08 => INIT_L_TH0_08,
      INIT_09 => INIT_L_TH0_09,
      INIT_0A => INIT_L_TH0_0A,
      INIT_0B => INIT_L_TH0_0B,
      INIT_0C => INIT_L_TH0_0C,
      INIT_0D => INIT_L_TH0_0D,
      INIT_0E => INIT_L_TH0_0E,
      INIT_0F => INIT_L_TH0_0F,
      INIT_10 => INIT_L_TH0_10,
      INIT_11 => INIT_L_TH0_11,
      INIT_12 => INIT_L_TH0_12,
      INIT_13 => INIT_L_TH0_13,
      INIT_14 => INIT_L_TH0_14,
      INIT_15 => INIT_L_TH0_15,
      INIT_16 => INIT_L_TH0_16,
      INIT_17 => INIT_L_TH0_17,
      INIT_18 => INIT_L_TH0_18,
      INIT_19 => INIT_L_TH0_19,
      INIT_1A => INIT_L_TH0_1A,
      INIT_1B => INIT_L_TH0_1B,
      INIT_1C => INIT_L_TH0_1C,
      INIT_1D => INIT_L_TH0_1D,
      INIT_1E => INIT_L_TH0_1E,
      INIT_1F => INIT_L_TH0_1F,
      INIT_20 => INIT_L_TH0_20,
      INIT_21 => INIT_L_TH0_21,
      INIT_22 => INIT_L_TH0_22,
      INIT_23 => INIT_L_TH0_23,
      INIT_24 => INIT_L_TH0_24,
      INIT_25 => INIT_L_TH0_25,
      INIT_26 => INIT_L_TH0_26,
      INIT_27 => INIT_L_TH0_27,
      INIT_28 => INIT_L_TH0_28,
      INIT_29 => INIT_L_TH0_29,
      INIT_2A => INIT_L_TH0_2A,
      INIT_2B => INIT_L_TH0_2B,
      INIT_2C => INIT_L_TH0_2C,
      INIT_2D => INIT_L_TH0_2D,
      INIT_2E => INIT_L_TH0_2E,
      INIT_2F => INIT_L_TH0_2F,
      INIT_30 => INIT_L_TH0_30,
      INIT_31 => INIT_L_TH0_31,
      INIT_32 => INIT_L_TH0_32,
      INIT_33 => INIT_L_TH0_33,
      INIT_34 => INIT_L_TH0_34,
      INIT_35 => INIT_L_TH0_35,
      INIT_36 => INIT_L_TH0_36,
      INIT_37 => INIT_L_TH0_37,
      INIT_38 => INIT_L_TH0_38,
      INIT_39 => INIT_L_TH0_39,
      INIT_3A => INIT_L_TH0_3A,
      INIT_3B => INIT_L_TH0_3B,
      INIT_3C => INIT_L_TH0_3C,
      INIT_3D => INIT_L_TH0_3D,
      INIT_3E => INIT_L_TH0_3E,
      INIT_3F => INIT_L_TH0_3F,
      INIT_40 => INIT_L_TH0_40,
      INIT_41 => INIT_L_TH0_41,
      INIT_42 => INIT_L_TH0_42,
      INIT_43 => INIT_L_TH0_43,
      INIT_44 => INIT_L_TH0_44,
      INIT_45 => INIT_L_TH0_45,
      INIT_46 => INIT_L_TH0_46,
      INIT_47 => INIT_L_TH0_47,
      INIT_48 => INIT_L_TH0_48,
      INIT_49 => INIT_L_TH0_49,
      INIT_4A => INIT_L_TH0_4A,
      INIT_4B => INIT_L_TH0_4B,
      INIT_4C => INIT_L_TH0_4C,
      INIT_4D => INIT_L_TH0_4D,
      INIT_4E => INIT_L_TH0_4E,
      INIT_4F => INIT_L_TH0_4F,
      INIT_50 => INIT_L_TH0_50,
      INIT_51 => INIT_L_TH0_51,
      INIT_52 => INIT_L_TH0_52,
      INIT_53 => INIT_L_TH0_53,
      INIT_54 => INIT_L_TH0_54,
      INIT_55 => INIT_L_TH0_55,
      INIT_56 => INIT_L_TH0_56,
      INIT_57 => INIT_L_TH0_57,
      INIT_58 => INIT_L_TH0_58,
      INIT_59 => INIT_L_TH0_59,
      INIT_5A => INIT_L_TH0_5A,
      INIT_5B => INIT_L_TH0_5B,
      INIT_5C => INIT_L_TH0_5C,
      INIT_5D => INIT_L_TH0_5D,
      INIT_5E => INIT_L_TH0_5E,
      INIT_5F => INIT_L_TH0_5F,
      INIT_60 => INIT_L_TH0_60,
      INIT_61 => INIT_L_TH0_61,
      INIT_62 => INIT_L_TH0_62,
      INIT_63 => INIT_L_TH0_63,
      INIT_64 => INIT_L_TH0_64,
      INIT_65 => INIT_L_TH0_65,
      INIT_66 => INIT_L_TH0_66,
      INIT_67 => INIT_L_TH0_67,
      INIT_68 => INIT_L_TH0_68,
      INIT_69 => INIT_L_TH0_69,
      INIT_6A => INIT_L_TH0_6A,
      INIT_6B => INIT_L_TH0_6B,
      INIT_6C => INIT_L_TH0_6C,
      INIT_6D => INIT_L_TH0_6D,
      INIT_6E => INIT_L_TH0_6E,
      INIT_6F => INIT_L_TH0_6F,
      INIT_70 => INIT_L_TH0_70,
      INIT_71 => INIT_L_TH0_71,
      INIT_72 => INIT_L_TH0_72,
      INIT_73 => INIT_L_TH0_73,
      INIT_74 => INIT_L_TH0_74,
      INIT_75 => INIT_L_TH0_75,
      INIT_76 => INIT_L_TH0_76,
      INIT_77 => INIT_L_TH0_77,
      INIT_78 => INIT_L_TH0_78,
      INIT_79 => INIT_L_TH0_79,
      INIT_7A => INIT_L_TH0_7A,
      INIT_7B => INIT_L_TH0_7B,
      INIT_7C => INIT_L_TH0_7C,
      INIT_7D => INIT_L_TH0_7D,
      INIT_7E => INIT_L_TH0_7E,
      INIT_7F => INIT_L_TH0_7F
   ) port map(
      ADDRARDADDR    => th0_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => th0_l_data_out_a(31 downto 0),
      DOPADOP        => th0_l_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );

   th0_address_a <= '1' & adcData(0)(23 downto 12) & "111";
   th0_data_out_a <= th0_h_data_out_a(7 downto 0) & th0_l_data_out_a(7 downto 0);
   outEnvData(0) <= std_logic_vector(resize(signed(th0_data_out_a), 32));



   th1_h_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_H_TH1_00,
      INIT_01 => INIT_H_TH1_01,
      INIT_02 => INIT_H_TH1_02,
      INIT_03 => INIT_H_TH1_03,
      INIT_04 => INIT_H_TH1_04,
      INIT_05 => INIT_H_TH1_05,
      INIT_06 => INIT_H_TH1_06,
      INIT_07 => INIT_H_TH1_07,
      INIT_08 => INIT_H_TH1_08,
      INIT_09 => INIT_H_TH1_09,
      INIT_0A => INIT_H_TH1_0A,
      INIT_0B => INIT_H_TH1_0B,
      INIT_0C => INIT_H_TH1_0C,
      INIT_0D => INIT_H_TH1_0D,
      INIT_0E => INIT_H_TH1_0E,
      INIT_0F => INIT_H_TH1_0F,
      INIT_10 => INIT_H_TH1_10,
      INIT_11 => INIT_H_TH1_11,
      INIT_12 => INIT_H_TH1_12,
      INIT_13 => INIT_H_TH1_13,
      INIT_14 => INIT_H_TH1_14,
      INIT_15 => INIT_H_TH1_15,
      INIT_16 => INIT_H_TH1_16,
      INIT_17 => INIT_H_TH1_17,
      INIT_18 => INIT_H_TH1_18,
      INIT_19 => INIT_H_TH1_19,
      INIT_1A => INIT_H_TH1_1A,
      INIT_1B => INIT_H_TH1_1B,
      INIT_1C => INIT_H_TH1_1C,
      INIT_1D => INIT_H_TH1_1D,
      INIT_1E => INIT_H_TH1_1E,
      INIT_1F => INIT_H_TH1_1F,
      INIT_20 => INIT_H_TH1_20,
      INIT_21 => INIT_H_TH1_21,
      INIT_22 => INIT_H_TH1_22,
      INIT_23 => INIT_H_TH1_23,
      INIT_24 => INIT_H_TH1_24,
      INIT_25 => INIT_H_TH1_25,
      INIT_26 => INIT_H_TH1_26,
      INIT_27 => INIT_H_TH1_27,
      INIT_28 => INIT_H_TH1_28,
      INIT_29 => INIT_H_TH1_29,
      INIT_2A => INIT_H_TH1_2A,
      INIT_2B => INIT_H_TH1_2B,
      INIT_2C => INIT_H_TH1_2C,
      INIT_2D => INIT_H_TH1_2D,
      INIT_2E => INIT_H_TH1_2E,
      INIT_2F => INIT_H_TH1_2F,
      INIT_30 => INIT_H_TH1_30,
      INIT_31 => INIT_H_TH1_31,
      INIT_32 => INIT_H_TH1_32,
      INIT_33 => INIT_H_TH1_33,
      INIT_34 => INIT_H_TH1_34,
      INIT_35 => INIT_H_TH1_35,
      INIT_36 => INIT_H_TH1_36,
      INIT_37 => INIT_H_TH1_37,
      INIT_38 => INIT_H_TH1_38,
      INIT_39 => INIT_H_TH1_39,
      INIT_3A => INIT_H_TH1_3A,
      INIT_3B => INIT_H_TH1_3B,
      INIT_3C => INIT_H_TH1_3C,
      INIT_3D => INIT_H_TH1_3D,
      INIT_3E => INIT_H_TH1_3E,
      INIT_3F => INIT_H_TH1_3F,
      INIT_40 => INIT_H_TH1_40,
      INIT_41 => INIT_H_TH1_41,
      INIT_42 => INIT_H_TH1_42,
      INIT_43 => INIT_H_TH1_43,
      INIT_44 => INIT_H_TH1_44,
      INIT_45 => INIT_H_TH1_45,
      INIT_46 => INIT_H_TH1_46,
      INIT_47 => INIT_H_TH1_47,
      INIT_48 => INIT_H_TH1_48,
      INIT_49 => INIT_H_TH1_49,
      INIT_4A => INIT_H_TH1_4A,
      INIT_4B => INIT_H_TH1_4B,
      INIT_4C => INIT_H_TH1_4C,
      INIT_4D => INIT_H_TH1_4D,
      INIT_4E => INIT_H_TH1_4E,
      INIT_4F => INIT_H_TH1_4F,
      INIT_50 => INIT_H_TH1_50,
      INIT_51 => INIT_H_TH1_51,
      INIT_52 => INIT_H_TH1_52,
      INIT_53 => INIT_H_TH1_53,
      INIT_54 => INIT_H_TH1_54,
      INIT_55 => INIT_H_TH1_55,
      INIT_56 => INIT_H_TH1_56,
      INIT_57 => INIT_H_TH1_57,
      INIT_58 => INIT_H_TH1_58,
      INIT_59 => INIT_H_TH1_59,
      INIT_5A => INIT_H_TH1_5A,
      INIT_5B => INIT_H_TH1_5B,
      INIT_5C => INIT_H_TH1_5C,
      INIT_5D => INIT_H_TH1_5D,
      INIT_5E => INIT_H_TH1_5E,
      INIT_5F => INIT_H_TH1_5F,
      INIT_60 => INIT_H_TH1_60,
      INIT_61 => INIT_H_TH1_61,
      INIT_62 => INIT_H_TH1_62,
      INIT_63 => INIT_H_TH1_63,
      INIT_64 => INIT_H_TH1_64,
      INIT_65 => INIT_H_TH1_65,
      INIT_66 => INIT_H_TH1_66,
      INIT_67 => INIT_H_TH1_67,
      INIT_68 => INIT_H_TH1_68,
      INIT_69 => INIT_H_TH1_69,
      INIT_6A => INIT_H_TH1_6A,
      INIT_6B => INIT_H_TH1_6B,
      INIT_6C => INIT_H_TH1_6C,
      INIT_6D => INIT_H_TH1_6D,
      INIT_6E => INIT_H_TH1_6E,
      INIT_6F => INIT_H_TH1_6F,
      INIT_70 => INIT_H_TH1_70,
      INIT_71 => INIT_H_TH1_71,
      INIT_72 => INIT_H_TH1_72,
      INIT_73 => INIT_H_TH1_73,
      INIT_74 => INIT_H_TH1_74,
      INIT_75 => INIT_H_TH1_75,
      INIT_76 => INIT_H_TH1_76,
      INIT_77 => INIT_H_TH1_77,
      INIT_78 => INIT_H_TH1_78,
      INIT_79 => INIT_H_TH1_79,
      INIT_7A => INIT_H_TH1_7A,
      INIT_7B => INIT_H_TH1_7B,
      INIT_7C => INIT_H_TH1_7C,
      INIT_7D => INIT_H_TH1_7D,
      INIT_7E => INIT_H_TH1_7E,
      INIT_7F => INIT_H_TH1_7F
   ) port map(
      ADDRARDADDR    => th1_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => th1_h_data_out_a(31 downto 0),
      DOPADOP        => th1_h_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );



   th1_l_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_L_TH1_00,
      INIT_01 => INIT_L_TH1_01,
      INIT_02 => INIT_L_TH1_02,
      INIT_03 => INIT_L_TH1_03,
      INIT_04 => INIT_L_TH1_04,
      INIT_05 => INIT_L_TH1_05,
      INIT_06 => INIT_L_TH1_06,
      INIT_07 => INIT_L_TH1_07,
      INIT_08 => INIT_L_TH1_08,
      INIT_09 => INIT_L_TH1_09,
      INIT_0A => INIT_L_TH1_0A,
      INIT_0B => INIT_L_TH1_0B,
      INIT_0C => INIT_L_TH1_0C,
      INIT_0D => INIT_L_TH1_0D,
      INIT_0E => INIT_L_TH1_0E,
      INIT_0F => INIT_L_TH1_0F,
      INIT_10 => INIT_L_TH1_10,
      INIT_11 => INIT_L_TH1_11,
      INIT_12 => INIT_L_TH1_12,
      INIT_13 => INIT_L_TH1_13,
      INIT_14 => INIT_L_TH1_14,
      INIT_15 => INIT_L_TH1_15,
      INIT_16 => INIT_L_TH1_16,
      INIT_17 => INIT_L_TH1_17,
      INIT_18 => INIT_L_TH1_18,
      INIT_19 => INIT_L_TH1_19,
      INIT_1A => INIT_L_TH1_1A,
      INIT_1B => INIT_L_TH1_1B,
      INIT_1C => INIT_L_TH1_1C,
      INIT_1D => INIT_L_TH1_1D,
      INIT_1E => INIT_L_TH1_1E,
      INIT_1F => INIT_L_TH1_1F,
      INIT_20 => INIT_L_TH1_20,
      INIT_21 => INIT_L_TH1_21,
      INIT_22 => INIT_L_TH1_22,
      INIT_23 => INIT_L_TH1_23,
      INIT_24 => INIT_L_TH1_24,
      INIT_25 => INIT_L_TH1_25,
      INIT_26 => INIT_L_TH1_26,
      INIT_27 => INIT_L_TH1_27,
      INIT_28 => INIT_L_TH1_28,
      INIT_29 => INIT_L_TH1_29,
      INIT_2A => INIT_L_TH1_2A,
      INIT_2B => INIT_L_TH1_2B,
      INIT_2C => INIT_L_TH1_2C,
      INIT_2D => INIT_L_TH1_2D,
      INIT_2E => INIT_L_TH1_2E,
      INIT_2F => INIT_L_TH1_2F,
      INIT_30 => INIT_L_TH1_30,
      INIT_31 => INIT_L_TH1_31,
      INIT_32 => INIT_L_TH1_32,
      INIT_33 => INIT_L_TH1_33,
      INIT_34 => INIT_L_TH1_34,
      INIT_35 => INIT_L_TH1_35,
      INIT_36 => INIT_L_TH1_36,
      INIT_37 => INIT_L_TH1_37,
      INIT_38 => INIT_L_TH1_38,
      INIT_39 => INIT_L_TH1_39,
      INIT_3A => INIT_L_TH1_3A,
      INIT_3B => INIT_L_TH1_3B,
      INIT_3C => INIT_L_TH1_3C,
      INIT_3D => INIT_L_TH1_3D,
      INIT_3E => INIT_L_TH1_3E,
      INIT_3F => INIT_L_TH1_3F,
      INIT_40 => INIT_L_TH1_40,
      INIT_41 => INIT_L_TH1_41,
      INIT_42 => INIT_L_TH1_42,
      INIT_43 => INIT_L_TH1_43,
      INIT_44 => INIT_L_TH1_44,
      INIT_45 => INIT_L_TH1_45,
      INIT_46 => INIT_L_TH1_46,
      INIT_47 => INIT_L_TH1_47,
      INIT_48 => INIT_L_TH1_48,
      INIT_49 => INIT_L_TH1_49,
      INIT_4A => INIT_L_TH1_4A,
      INIT_4B => INIT_L_TH1_4B,
      INIT_4C => INIT_L_TH1_4C,
      INIT_4D => INIT_L_TH1_4D,
      INIT_4E => INIT_L_TH1_4E,
      INIT_4F => INIT_L_TH1_4F,
      INIT_50 => INIT_L_TH1_50,
      INIT_51 => INIT_L_TH1_51,
      INIT_52 => INIT_L_TH1_52,
      INIT_53 => INIT_L_TH1_53,
      INIT_54 => INIT_L_TH1_54,
      INIT_55 => INIT_L_TH1_55,
      INIT_56 => INIT_L_TH1_56,
      INIT_57 => INIT_L_TH1_57,
      INIT_58 => INIT_L_TH1_58,
      INIT_59 => INIT_L_TH1_59,
      INIT_5A => INIT_L_TH1_5A,
      INIT_5B => INIT_L_TH1_5B,
      INIT_5C => INIT_L_TH1_5C,
      INIT_5D => INIT_L_TH1_5D,
      INIT_5E => INIT_L_TH1_5E,
      INIT_5F => INIT_L_TH1_5F,
      INIT_60 => INIT_L_TH1_60,
      INIT_61 => INIT_L_TH1_61,
      INIT_62 => INIT_L_TH1_62,
      INIT_63 => INIT_L_TH1_63,
      INIT_64 => INIT_L_TH1_64,
      INIT_65 => INIT_L_TH1_65,
      INIT_66 => INIT_L_TH1_66,
      INIT_67 => INIT_L_TH1_67,
      INIT_68 => INIT_L_TH1_68,
      INIT_69 => INIT_L_TH1_69,
      INIT_6A => INIT_L_TH1_6A,
      INIT_6B => INIT_L_TH1_6B,
      INIT_6C => INIT_L_TH1_6C,
      INIT_6D => INIT_L_TH1_6D,
      INIT_6E => INIT_L_TH1_6E,
      INIT_6F => INIT_L_TH1_6F,
      INIT_70 => INIT_L_TH1_70,
      INIT_71 => INIT_L_TH1_71,
      INIT_72 => INIT_L_TH1_72,
      INIT_73 => INIT_L_TH1_73,
      INIT_74 => INIT_L_TH1_74,
      INIT_75 => INIT_L_TH1_75,
      INIT_76 => INIT_L_TH1_76,
      INIT_77 => INIT_L_TH1_77,
      INIT_78 => INIT_L_TH1_78,
      INIT_79 => INIT_L_TH1_79,
      INIT_7A => INIT_L_TH1_7A,
      INIT_7B => INIT_L_TH1_7B,
      INIT_7C => INIT_L_TH1_7C,
      INIT_7D => INIT_L_TH1_7D,
      INIT_7E => INIT_L_TH1_7E,
      INIT_7F => INIT_L_TH1_7F
   ) port map(
      ADDRARDADDR    => th1_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => th1_l_data_out_a(31 downto 0),
      DOPADOP        => th1_l_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );

   th1_address_a <= '1' & adcData(1)(23 downto 12) & "111";
   th1_data_out_a <= th1_h_data_out_a(7 downto 0) & th1_l_data_out_a(7 downto 0);
   outEnvData(1) <= std_logic_vector(resize(signed(th1_data_out_a), 32));


   hum_h_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_H_HUM_00,
      INIT_01 => INIT_H_HUM_01,
      INIT_02 => INIT_H_HUM_02,
      INIT_03 => INIT_H_HUM_03,
      INIT_04 => INIT_H_HUM_04,
      INIT_05 => INIT_H_HUM_05,
      INIT_06 => INIT_H_HUM_06,
      INIT_07 => INIT_H_HUM_07,
      INIT_08 => INIT_H_HUM_08,
      INIT_09 => INIT_H_HUM_09,
      INIT_0A => INIT_H_HUM_0A,
      INIT_0B => INIT_H_HUM_0B,
      INIT_0C => INIT_H_HUM_0C,
      INIT_0D => INIT_H_HUM_0D,
      INIT_0E => INIT_H_HUM_0E,
      INIT_0F => INIT_H_HUM_0F,
      INIT_10 => INIT_H_HUM_10,
      INIT_11 => INIT_H_HUM_11,
      INIT_12 => INIT_H_HUM_12,
      INIT_13 => INIT_H_HUM_13,
      INIT_14 => INIT_H_HUM_14,
      INIT_15 => INIT_H_HUM_15,
      INIT_16 => INIT_H_HUM_16,
      INIT_17 => INIT_H_HUM_17,
      INIT_18 => INIT_H_HUM_18,
      INIT_19 => INIT_H_HUM_19,
      INIT_1A => INIT_H_HUM_1A,
      INIT_1B => INIT_H_HUM_1B,
      INIT_1C => INIT_H_HUM_1C,
      INIT_1D => INIT_H_HUM_1D,
      INIT_1E => INIT_H_HUM_1E,
      INIT_1F => INIT_H_HUM_1F,
      INIT_20 => INIT_H_HUM_20,
      INIT_21 => INIT_H_HUM_21,
      INIT_22 => INIT_H_HUM_22,
      INIT_23 => INIT_H_HUM_23,
      INIT_24 => INIT_H_HUM_24,
      INIT_25 => INIT_H_HUM_25,
      INIT_26 => INIT_H_HUM_26,
      INIT_27 => INIT_H_HUM_27,
      INIT_28 => INIT_H_HUM_28,
      INIT_29 => INIT_H_HUM_29,
      INIT_2A => INIT_H_HUM_2A,
      INIT_2B => INIT_H_HUM_2B,
      INIT_2C => INIT_H_HUM_2C,
      INIT_2D => INIT_H_HUM_2D,
      INIT_2E => INIT_H_HUM_2E,
      INIT_2F => INIT_H_HUM_2F,
      INIT_30 => INIT_H_HUM_30,
      INIT_31 => INIT_H_HUM_31,
      INIT_32 => INIT_H_HUM_32,
      INIT_33 => INIT_H_HUM_33,
      INIT_34 => INIT_H_HUM_34,
      INIT_35 => INIT_H_HUM_35,
      INIT_36 => INIT_H_HUM_36,
      INIT_37 => INIT_H_HUM_37,
      INIT_38 => INIT_H_HUM_38,
      INIT_39 => INIT_H_HUM_39,
      INIT_3A => INIT_H_HUM_3A,
      INIT_3B => INIT_H_HUM_3B,
      INIT_3C => INIT_H_HUM_3C,
      INIT_3D => INIT_H_HUM_3D,
      INIT_3E => INIT_H_HUM_3E,
      INIT_3F => INIT_H_HUM_3F,
      INIT_40 => INIT_H_HUM_40,
      INIT_41 => INIT_H_HUM_41,
      INIT_42 => INIT_H_HUM_42,
      INIT_43 => INIT_H_HUM_43,
      INIT_44 => INIT_H_HUM_44,
      INIT_45 => INIT_H_HUM_45,
      INIT_46 => INIT_H_HUM_46,
      INIT_47 => INIT_H_HUM_47,
      INIT_48 => INIT_H_HUM_48,
      INIT_49 => INIT_H_HUM_49,
      INIT_4A => INIT_H_HUM_4A,
      INIT_4B => INIT_H_HUM_4B,
      INIT_4C => INIT_H_HUM_4C,
      INIT_4D => INIT_H_HUM_4D,
      INIT_4E => INIT_H_HUM_4E,
      INIT_4F => INIT_H_HUM_4F,
      INIT_50 => INIT_H_HUM_50,
      INIT_51 => INIT_H_HUM_51,
      INIT_52 => INIT_H_HUM_52,
      INIT_53 => INIT_H_HUM_53,
      INIT_54 => INIT_H_HUM_54,
      INIT_55 => INIT_H_HUM_55,
      INIT_56 => INIT_H_HUM_56,
      INIT_57 => INIT_H_HUM_57,
      INIT_58 => INIT_H_HUM_58,
      INIT_59 => INIT_H_HUM_59,
      INIT_5A => INIT_H_HUM_5A,
      INIT_5B => INIT_H_HUM_5B,
      INIT_5C => INIT_H_HUM_5C,
      INIT_5D => INIT_H_HUM_5D,
      INIT_5E => INIT_H_HUM_5E,
      INIT_5F => INIT_H_HUM_5F,
      INIT_60 => INIT_H_HUM_60,
      INIT_61 => INIT_H_HUM_61,
      INIT_62 => INIT_H_HUM_62,
      INIT_63 => INIT_H_HUM_63,
      INIT_64 => INIT_H_HUM_64,
      INIT_65 => INIT_H_HUM_65,
      INIT_66 => INIT_H_HUM_66,
      INIT_67 => INIT_H_HUM_67,
      INIT_68 => INIT_H_HUM_68,
      INIT_69 => INIT_H_HUM_69,
      INIT_6A => INIT_H_HUM_6A,
      INIT_6B => INIT_H_HUM_6B,
      INIT_6C => INIT_H_HUM_6C,
      INIT_6D => INIT_H_HUM_6D,
      INIT_6E => INIT_H_HUM_6E,
      INIT_6F => INIT_H_HUM_6F,
      INIT_70 => INIT_H_HUM_70,
      INIT_71 => INIT_H_HUM_71,
      INIT_72 => INIT_H_HUM_72,
      INIT_73 => INIT_H_HUM_73,
      INIT_74 => INIT_H_HUM_74,
      INIT_75 => INIT_H_HUM_75,
      INIT_76 => INIT_H_HUM_76,
      INIT_77 => INIT_H_HUM_77,
      INIT_78 => INIT_H_HUM_78,
      INIT_79 => INIT_H_HUM_79,
      INIT_7A => INIT_H_HUM_7A,
      INIT_7B => INIT_H_HUM_7B,
      INIT_7C => INIT_H_HUM_7C,
      INIT_7D => INIT_H_HUM_7D,
      INIT_7E => INIT_H_HUM_7E,
      INIT_7F => INIT_H_HUM_7F
   ) port map(
      ADDRARDADDR    => hum_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => hum_h_data_out_a(31 downto 0),
      DOPADOP        => hum_h_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );



   hum_l_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_L_HUM_00,
      INIT_01 => INIT_L_HUM_01,
      INIT_02 => INIT_L_HUM_02,
      INIT_03 => INIT_L_HUM_03,
      INIT_04 => INIT_L_HUM_04,
      INIT_05 => INIT_L_HUM_05,
      INIT_06 => INIT_L_HUM_06,
      INIT_07 => INIT_L_HUM_07,
      INIT_08 => INIT_L_HUM_08,
      INIT_09 => INIT_L_HUM_09,
      INIT_0A => INIT_L_HUM_0A,
      INIT_0B => INIT_L_HUM_0B,
      INIT_0C => INIT_L_HUM_0C,
      INIT_0D => INIT_L_HUM_0D,
      INIT_0E => INIT_L_HUM_0E,
      INIT_0F => INIT_L_HUM_0F,
      INIT_10 => INIT_L_HUM_10,
      INIT_11 => INIT_L_HUM_11,
      INIT_12 => INIT_L_HUM_12,
      INIT_13 => INIT_L_HUM_13,
      INIT_14 => INIT_L_HUM_14,
      INIT_15 => INIT_L_HUM_15,
      INIT_16 => INIT_L_HUM_16,
      INIT_17 => INIT_L_HUM_17,
      INIT_18 => INIT_L_HUM_18,
      INIT_19 => INIT_L_HUM_19,
      INIT_1A => INIT_L_HUM_1A,
      INIT_1B => INIT_L_HUM_1B,
      INIT_1C => INIT_L_HUM_1C,
      INIT_1D => INIT_L_HUM_1D,
      INIT_1E => INIT_L_HUM_1E,
      INIT_1F => INIT_L_HUM_1F,
      INIT_20 => INIT_L_HUM_20,
      INIT_21 => INIT_L_HUM_21,
      INIT_22 => INIT_L_HUM_22,
      INIT_23 => INIT_L_HUM_23,
      INIT_24 => INIT_L_HUM_24,
      INIT_25 => INIT_L_HUM_25,
      INIT_26 => INIT_L_HUM_26,
      INIT_27 => INIT_L_HUM_27,
      INIT_28 => INIT_L_HUM_28,
      INIT_29 => INIT_L_HUM_29,
      INIT_2A => INIT_L_HUM_2A,
      INIT_2B => INIT_L_HUM_2B,
      INIT_2C => INIT_L_HUM_2C,
      INIT_2D => INIT_L_HUM_2D,
      INIT_2E => INIT_L_HUM_2E,
      INIT_2F => INIT_L_HUM_2F,
      INIT_30 => INIT_L_HUM_30,
      INIT_31 => INIT_L_HUM_31,
      INIT_32 => INIT_L_HUM_32,
      INIT_33 => INIT_L_HUM_33,
      INIT_34 => INIT_L_HUM_34,
      INIT_35 => INIT_L_HUM_35,
      INIT_36 => INIT_L_HUM_36,
      INIT_37 => INIT_L_HUM_37,
      INIT_38 => INIT_L_HUM_38,
      INIT_39 => INIT_L_HUM_39,
      INIT_3A => INIT_L_HUM_3A,
      INIT_3B => INIT_L_HUM_3B,
      INIT_3C => INIT_L_HUM_3C,
      INIT_3D => INIT_L_HUM_3D,
      INIT_3E => INIT_L_HUM_3E,
      INIT_3F => INIT_L_HUM_3F,
      INIT_40 => INIT_L_HUM_40,
      INIT_41 => INIT_L_HUM_41,
      INIT_42 => INIT_L_HUM_42,
      INIT_43 => INIT_L_HUM_43,
      INIT_44 => INIT_L_HUM_44,
      INIT_45 => INIT_L_HUM_45,
      INIT_46 => INIT_L_HUM_46,
      INIT_47 => INIT_L_HUM_47,
      INIT_48 => INIT_L_HUM_48,
      INIT_49 => INIT_L_HUM_49,
      INIT_4A => INIT_L_HUM_4A,
      INIT_4B => INIT_L_HUM_4B,
      INIT_4C => INIT_L_HUM_4C,
      INIT_4D => INIT_L_HUM_4D,
      INIT_4E => INIT_L_HUM_4E,
      INIT_4F => INIT_L_HUM_4F,
      INIT_50 => INIT_L_HUM_50,
      INIT_51 => INIT_L_HUM_51,
      INIT_52 => INIT_L_HUM_52,
      INIT_53 => INIT_L_HUM_53,
      INIT_54 => INIT_L_HUM_54,
      INIT_55 => INIT_L_HUM_55,
      INIT_56 => INIT_L_HUM_56,
      INIT_57 => INIT_L_HUM_57,
      INIT_58 => INIT_L_HUM_58,
      INIT_59 => INIT_L_HUM_59,
      INIT_5A => INIT_L_HUM_5A,
      INIT_5B => INIT_L_HUM_5B,
      INIT_5C => INIT_L_HUM_5C,
      INIT_5D => INIT_L_HUM_5D,
      INIT_5E => INIT_L_HUM_5E,
      INIT_5F => INIT_L_HUM_5F,
      INIT_60 => INIT_L_HUM_60,
      INIT_61 => INIT_L_HUM_61,
      INIT_62 => INIT_L_HUM_62,
      INIT_63 => INIT_L_HUM_63,
      INIT_64 => INIT_L_HUM_64,
      INIT_65 => INIT_L_HUM_65,
      INIT_66 => INIT_L_HUM_66,
      INIT_67 => INIT_L_HUM_67,
      INIT_68 => INIT_L_HUM_68,
      INIT_69 => INIT_L_HUM_69,
      INIT_6A => INIT_L_HUM_6A,
      INIT_6B => INIT_L_HUM_6B,
      INIT_6C => INIT_L_HUM_6C,
      INIT_6D => INIT_L_HUM_6D,
      INIT_6E => INIT_L_HUM_6E,
      INIT_6F => INIT_L_HUM_6F,
      INIT_70 => INIT_L_HUM_70,
      INIT_71 => INIT_L_HUM_71,
      INIT_72 => INIT_L_HUM_72,
      INIT_73 => INIT_L_HUM_73,
      INIT_74 => INIT_L_HUM_74,
      INIT_75 => INIT_L_HUM_75,
      INIT_76 => INIT_L_HUM_76,
      INIT_77 => INIT_L_HUM_77,
      INIT_78 => INIT_L_HUM_78,
      INIT_79 => INIT_L_HUM_79,
      INIT_7A => INIT_L_HUM_7A,
      INIT_7B => INIT_L_HUM_7B,
      INIT_7C => INIT_L_HUM_7C,
      INIT_7D => INIT_L_HUM_7D,
      INIT_7E => INIT_L_HUM_7E,
      INIT_7F => INIT_L_HUM_7F
   ) port map(
      ADDRARDADDR    => hum_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => hum_l_data_out_a(31 downto 0),
      DOPADOP        => hum_l_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );

   hum_address_a <= '1' & adcData(2)(23 downto 12) & "111";
   hum_data_out_a <= hum_h_data_out_a(7 downto 0) & hum_l_data_out_a(7 downto 0);
   outEnvData(2) <= std_logic_vector(resize(signed(hum_data_out_a), 32));

   iana_h_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_H_IANA_00,
      INIT_01 => INIT_H_IANA_01,
      INIT_02 => INIT_H_IANA_02,
      INIT_03 => INIT_H_IANA_03,
      INIT_04 => INIT_H_IANA_04,
      INIT_05 => INIT_H_IANA_05,
      INIT_06 => INIT_H_IANA_06,
      INIT_07 => INIT_H_IANA_07,
      INIT_08 => INIT_H_IANA_08,
      INIT_09 => INIT_H_IANA_09,
      INIT_0A => INIT_H_IANA_0A,
      INIT_0B => INIT_H_IANA_0B,
      INIT_0C => INIT_H_IANA_0C,
      INIT_0D => INIT_H_IANA_0D,
      INIT_0E => INIT_H_IANA_0E,
      INIT_0F => INIT_H_IANA_0F,
      INIT_10 => INIT_H_IANA_10,
      INIT_11 => INIT_H_IANA_11,
      INIT_12 => INIT_H_IANA_12,
      INIT_13 => INIT_H_IANA_13,
      INIT_14 => INIT_H_IANA_14,
      INIT_15 => INIT_H_IANA_15,
      INIT_16 => INIT_H_IANA_16,
      INIT_17 => INIT_H_IANA_17,
      INIT_18 => INIT_H_IANA_18,
      INIT_19 => INIT_H_IANA_19,
      INIT_1A => INIT_H_IANA_1A,
      INIT_1B => INIT_H_IANA_1B,
      INIT_1C => INIT_H_IANA_1C,
      INIT_1D => INIT_H_IANA_1D,
      INIT_1E => INIT_H_IANA_1E,
      INIT_1F => INIT_H_IANA_1F,
      INIT_20 => INIT_H_IANA_20,
      INIT_21 => INIT_H_IANA_21,
      INIT_22 => INIT_H_IANA_22,
      INIT_23 => INIT_H_IANA_23,
      INIT_24 => INIT_H_IANA_24,
      INIT_25 => INIT_H_IANA_25,
      INIT_26 => INIT_H_IANA_26,
      INIT_27 => INIT_H_IANA_27,
      INIT_28 => INIT_H_IANA_28,
      INIT_29 => INIT_H_IANA_29,
      INIT_2A => INIT_H_IANA_2A,
      INIT_2B => INIT_H_IANA_2B,
      INIT_2C => INIT_H_IANA_2C,
      INIT_2D => INIT_H_IANA_2D,
      INIT_2E => INIT_H_IANA_2E,
      INIT_2F => INIT_H_IANA_2F,
      INIT_30 => INIT_H_IANA_30,
      INIT_31 => INIT_H_IANA_31,
      INIT_32 => INIT_H_IANA_32,
      INIT_33 => INIT_H_IANA_33,
      INIT_34 => INIT_H_IANA_34,
      INIT_35 => INIT_H_IANA_35,
      INIT_36 => INIT_H_IANA_36,
      INIT_37 => INIT_H_IANA_37,
      INIT_38 => INIT_H_IANA_38,
      INIT_39 => INIT_H_IANA_39,
      INIT_3A => INIT_H_IANA_3A,
      INIT_3B => INIT_H_IANA_3B,
      INIT_3C => INIT_H_IANA_3C,
      INIT_3D => INIT_H_IANA_3D,
      INIT_3E => INIT_H_IANA_3E,
      INIT_3F => INIT_H_IANA_3F,
      INIT_40 => INIT_H_IANA_40,
      INIT_41 => INIT_H_IANA_41,
      INIT_42 => INIT_H_IANA_42,
      INIT_43 => INIT_H_IANA_43,
      INIT_44 => INIT_H_IANA_44,
      INIT_45 => INIT_H_IANA_45,
      INIT_46 => INIT_H_IANA_46,
      INIT_47 => INIT_H_IANA_47,
      INIT_48 => INIT_H_IANA_48,
      INIT_49 => INIT_H_IANA_49,
      INIT_4A => INIT_H_IANA_4A,
      INIT_4B => INIT_H_IANA_4B,
      INIT_4C => INIT_H_IANA_4C,
      INIT_4D => INIT_H_IANA_4D,
      INIT_4E => INIT_H_IANA_4E,
      INIT_4F => INIT_H_IANA_4F,
      INIT_50 => INIT_H_IANA_50,
      INIT_51 => INIT_H_IANA_51,
      INIT_52 => INIT_H_IANA_52,
      INIT_53 => INIT_H_IANA_53,
      INIT_54 => INIT_H_IANA_54,
      INIT_55 => INIT_H_IANA_55,
      INIT_56 => INIT_H_IANA_56,
      INIT_57 => INIT_H_IANA_57,
      INIT_58 => INIT_H_IANA_58,
      INIT_59 => INIT_H_IANA_59,
      INIT_5A => INIT_H_IANA_5A,
      INIT_5B => INIT_H_IANA_5B,
      INIT_5C => INIT_H_IANA_5C,
      INIT_5D => INIT_H_IANA_5D,
      INIT_5E => INIT_H_IANA_5E,
      INIT_5F => INIT_H_IANA_5F,
      INIT_60 => INIT_H_IANA_60,
      INIT_61 => INIT_H_IANA_61,
      INIT_62 => INIT_H_IANA_62,
      INIT_63 => INIT_H_IANA_63,
      INIT_64 => INIT_H_IANA_64,
      INIT_65 => INIT_H_IANA_65,
      INIT_66 => INIT_H_IANA_66,
      INIT_67 => INIT_H_IANA_67,
      INIT_68 => INIT_H_IANA_68,
      INIT_69 => INIT_H_IANA_69,
      INIT_6A => INIT_H_IANA_6A,
      INIT_6B => INIT_H_IANA_6B,
      INIT_6C => INIT_H_IANA_6C,
      INIT_6D => INIT_H_IANA_6D,
      INIT_6E => INIT_H_IANA_6E,
      INIT_6F => INIT_H_IANA_6F,
      INIT_70 => INIT_H_IANA_70,
      INIT_71 => INIT_H_IANA_71,
      INIT_72 => INIT_H_IANA_72,
      INIT_73 => INIT_H_IANA_73,
      INIT_74 => INIT_H_IANA_74,
      INIT_75 => INIT_H_IANA_75,
      INIT_76 => INIT_H_IANA_76,
      INIT_77 => INIT_H_IANA_77,
      INIT_78 => INIT_H_IANA_78,
      INIT_79 => INIT_H_IANA_79,
      INIT_7A => INIT_H_IANA_7A,
      INIT_7B => INIT_H_IANA_7B,
      INIT_7C => INIT_H_IANA_7C,
      INIT_7D => INIT_H_IANA_7D,
      INIT_7E => INIT_H_IANA_7E,
      INIT_7F => INIT_H_IANA_7F
   ) port map(
      ADDRARDADDR    => iana_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => iana_h_data_out_a(31 downto 0),
      DOPADOP        => iana_h_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );



   iana_l_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_L_IANA_00,
      INIT_01 => INIT_L_IANA_01,
      INIT_02 => INIT_L_IANA_02,
      INIT_03 => INIT_L_IANA_03,
      INIT_04 => INIT_L_IANA_04,
      INIT_05 => INIT_L_IANA_05,
      INIT_06 => INIT_L_IANA_06,
      INIT_07 => INIT_L_IANA_07,
      INIT_08 => INIT_L_IANA_08,
      INIT_09 => INIT_L_IANA_09,
      INIT_0A => INIT_L_IANA_0A,
      INIT_0B => INIT_L_IANA_0B,
      INIT_0C => INIT_L_IANA_0C,
      INIT_0D => INIT_L_IANA_0D,
      INIT_0E => INIT_L_IANA_0E,
      INIT_0F => INIT_L_IANA_0F,
      INIT_10 => INIT_L_IANA_10,
      INIT_11 => INIT_L_IANA_11,
      INIT_12 => INIT_L_IANA_12,
      INIT_13 => INIT_L_IANA_13,
      INIT_14 => INIT_L_IANA_14,
      INIT_15 => INIT_L_IANA_15,
      INIT_16 => INIT_L_IANA_16,
      INIT_17 => INIT_L_IANA_17,
      INIT_18 => INIT_L_IANA_18,
      INIT_19 => INIT_L_IANA_19,
      INIT_1A => INIT_L_IANA_1A,
      INIT_1B => INIT_L_IANA_1B,
      INIT_1C => INIT_L_IANA_1C,
      INIT_1D => INIT_L_IANA_1D,
      INIT_1E => INIT_L_IANA_1E,
      INIT_1F => INIT_L_IANA_1F,
      INIT_20 => INIT_L_IANA_20,
      INIT_21 => INIT_L_IANA_21,
      INIT_22 => INIT_L_IANA_22,
      INIT_23 => INIT_L_IANA_23,
      INIT_24 => INIT_L_IANA_24,
      INIT_25 => INIT_L_IANA_25,
      INIT_26 => INIT_L_IANA_26,
      INIT_27 => INIT_L_IANA_27,
      INIT_28 => INIT_L_IANA_28,
      INIT_29 => INIT_L_IANA_29,
      INIT_2A => INIT_L_IANA_2A,
      INIT_2B => INIT_L_IANA_2B,
      INIT_2C => INIT_L_IANA_2C,
      INIT_2D => INIT_L_IANA_2D,
      INIT_2E => INIT_L_IANA_2E,
      INIT_2F => INIT_L_IANA_2F,
      INIT_30 => INIT_L_IANA_30,
      INIT_31 => INIT_L_IANA_31,
      INIT_32 => INIT_L_IANA_32,
      INIT_33 => INIT_L_IANA_33,
      INIT_34 => INIT_L_IANA_34,
      INIT_35 => INIT_L_IANA_35,
      INIT_36 => INIT_L_IANA_36,
      INIT_37 => INIT_L_IANA_37,
      INIT_38 => INIT_L_IANA_38,
      INIT_39 => INIT_L_IANA_39,
      INIT_3A => INIT_L_IANA_3A,
      INIT_3B => INIT_L_IANA_3B,
      INIT_3C => INIT_L_IANA_3C,
      INIT_3D => INIT_L_IANA_3D,
      INIT_3E => INIT_L_IANA_3E,
      INIT_3F => INIT_L_IANA_3F,
      INIT_40 => INIT_L_IANA_40,
      INIT_41 => INIT_L_IANA_41,
      INIT_42 => INIT_L_IANA_42,
      INIT_43 => INIT_L_IANA_43,
      INIT_44 => INIT_L_IANA_44,
      INIT_45 => INIT_L_IANA_45,
      INIT_46 => INIT_L_IANA_46,
      INIT_47 => INIT_L_IANA_47,
      INIT_48 => INIT_L_IANA_48,
      INIT_49 => INIT_L_IANA_49,
      INIT_4A => INIT_L_IANA_4A,
      INIT_4B => INIT_L_IANA_4B,
      INIT_4C => INIT_L_IANA_4C,
      INIT_4D => INIT_L_IANA_4D,
      INIT_4E => INIT_L_IANA_4E,
      INIT_4F => INIT_L_IANA_4F,
      INIT_50 => INIT_L_IANA_50,
      INIT_51 => INIT_L_IANA_51,
      INIT_52 => INIT_L_IANA_52,
      INIT_53 => INIT_L_IANA_53,
      INIT_54 => INIT_L_IANA_54,
      INIT_55 => INIT_L_IANA_55,
      INIT_56 => INIT_L_IANA_56,
      INIT_57 => INIT_L_IANA_57,
      INIT_58 => INIT_L_IANA_58,
      INIT_59 => INIT_L_IANA_59,
      INIT_5A => INIT_L_IANA_5A,
      INIT_5B => INIT_L_IANA_5B,
      INIT_5C => INIT_L_IANA_5C,
      INIT_5D => INIT_L_IANA_5D,
      INIT_5E => INIT_L_IANA_5E,
      INIT_5F => INIT_L_IANA_5F,
      INIT_60 => INIT_L_IANA_60,
      INIT_61 => INIT_L_IANA_61,
      INIT_62 => INIT_L_IANA_62,
      INIT_63 => INIT_L_IANA_63,
      INIT_64 => INIT_L_IANA_64,
      INIT_65 => INIT_L_IANA_65,
      INIT_66 => INIT_L_IANA_66,
      INIT_67 => INIT_L_IANA_67,
      INIT_68 => INIT_L_IANA_68,
      INIT_69 => INIT_L_IANA_69,
      INIT_6A => INIT_L_IANA_6A,
      INIT_6B => INIT_L_IANA_6B,
      INIT_6C => INIT_L_IANA_6C,
      INIT_6D => INIT_L_IANA_6D,
      INIT_6E => INIT_L_IANA_6E,
      INIT_6F => INIT_L_IANA_6F,
      INIT_70 => INIT_L_IANA_70,
      INIT_71 => INIT_L_IANA_71,
      INIT_72 => INIT_L_IANA_72,
      INIT_73 => INIT_L_IANA_73,
      INIT_74 => INIT_L_IANA_74,
      INIT_75 => INIT_L_IANA_75,
      INIT_76 => INIT_L_IANA_76,
      INIT_77 => INIT_L_IANA_77,
      INIT_78 => INIT_L_IANA_78,
      INIT_79 => INIT_L_IANA_79,
      INIT_7A => INIT_L_IANA_7A,
      INIT_7B => INIT_L_IANA_7B,
      INIT_7C => INIT_L_IANA_7C,
      INIT_7D => INIT_L_IANA_7D,
      INIT_7E => INIT_L_IANA_7E,
      INIT_7F => INIT_L_IANA_7F
   ) port map(
      ADDRARDADDR    => iana_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => iana_l_data_out_a(31 downto 0),
      DOPADOP        => iana_l_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );

   iana_address_a <= '1' & adcData(3)(23 downto 12) & "111";
   outEnvData(3) <= x"0000" & iana_h_data_out_a(7 downto 0) & iana_l_data_out_a(7 downto 0);


   idig_h_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_H_IDIG_00,
      INIT_01 => INIT_H_IDIG_01,
      INIT_02 => INIT_H_IDIG_02,
      INIT_03 => INIT_H_IDIG_03,
      INIT_04 => INIT_H_IDIG_04,
      INIT_05 => INIT_H_IDIG_05,
      INIT_06 => INIT_H_IDIG_06,
      INIT_07 => INIT_H_IDIG_07,
      INIT_08 => INIT_H_IDIG_08,
      INIT_09 => INIT_H_IDIG_09,
      INIT_0A => INIT_H_IDIG_0A,
      INIT_0B => INIT_H_IDIG_0B,
      INIT_0C => INIT_H_IDIG_0C,
      INIT_0D => INIT_H_IDIG_0D,
      INIT_0E => INIT_H_IDIG_0E,
      INIT_0F => INIT_H_IDIG_0F,
      INIT_10 => INIT_H_IDIG_10,
      INIT_11 => INIT_H_IDIG_11,
      INIT_12 => INIT_H_IDIG_12,
      INIT_13 => INIT_H_IDIG_13,
      INIT_14 => INIT_H_IDIG_14,
      INIT_15 => INIT_H_IDIG_15,
      INIT_16 => INIT_H_IDIG_16,
      INIT_17 => INIT_H_IDIG_17,
      INIT_18 => INIT_H_IDIG_18,
      INIT_19 => INIT_H_IDIG_19,
      INIT_1A => INIT_H_IDIG_1A,
      INIT_1B => INIT_H_IDIG_1B,
      INIT_1C => INIT_H_IDIG_1C,
      INIT_1D => INIT_H_IDIG_1D,
      INIT_1E => INIT_H_IDIG_1E,
      INIT_1F => INIT_H_IDIG_1F,
      INIT_20 => INIT_H_IDIG_20,
      INIT_21 => INIT_H_IDIG_21,
      INIT_22 => INIT_H_IDIG_22,
      INIT_23 => INIT_H_IDIG_23,
      INIT_24 => INIT_H_IDIG_24,
      INIT_25 => INIT_H_IDIG_25,
      INIT_26 => INIT_H_IDIG_26,
      INIT_27 => INIT_H_IDIG_27,
      INIT_28 => INIT_H_IDIG_28,
      INIT_29 => INIT_H_IDIG_29,
      INIT_2A => INIT_H_IDIG_2A,
      INIT_2B => INIT_H_IDIG_2B,
      INIT_2C => INIT_H_IDIG_2C,
      INIT_2D => INIT_H_IDIG_2D,
      INIT_2E => INIT_H_IDIG_2E,
      INIT_2F => INIT_H_IDIG_2F,
      INIT_30 => INIT_H_IDIG_30,
      INIT_31 => INIT_H_IDIG_31,
      INIT_32 => INIT_H_IDIG_32,
      INIT_33 => INIT_H_IDIG_33,
      INIT_34 => INIT_H_IDIG_34,
      INIT_35 => INIT_H_IDIG_35,
      INIT_36 => INIT_H_IDIG_36,
      INIT_37 => INIT_H_IDIG_37,
      INIT_38 => INIT_H_IDIG_38,
      INIT_39 => INIT_H_IDIG_39,
      INIT_3A => INIT_H_IDIG_3A,
      INIT_3B => INIT_H_IDIG_3B,
      INIT_3C => INIT_H_IDIG_3C,
      INIT_3D => INIT_H_IDIG_3D,
      INIT_3E => INIT_H_IDIG_3E,
      INIT_3F => INIT_H_IDIG_3F,
      INIT_40 => INIT_H_IDIG_40,
      INIT_41 => INIT_H_IDIG_41,
      INIT_42 => INIT_H_IDIG_42,
      INIT_43 => INIT_H_IDIG_43,
      INIT_44 => INIT_H_IDIG_44,
      INIT_45 => INIT_H_IDIG_45,
      INIT_46 => INIT_H_IDIG_46,
      INIT_47 => INIT_H_IDIG_47,
      INIT_48 => INIT_H_IDIG_48,
      INIT_49 => INIT_H_IDIG_49,
      INIT_4A => INIT_H_IDIG_4A,
      INIT_4B => INIT_H_IDIG_4B,
      INIT_4C => INIT_H_IDIG_4C,
      INIT_4D => INIT_H_IDIG_4D,
      INIT_4E => INIT_H_IDIG_4E,
      INIT_4F => INIT_H_IDIG_4F,
      INIT_50 => INIT_H_IDIG_50,
      INIT_51 => INIT_H_IDIG_51,
      INIT_52 => INIT_H_IDIG_52,
      INIT_53 => INIT_H_IDIG_53,
      INIT_54 => INIT_H_IDIG_54,
      INIT_55 => INIT_H_IDIG_55,
      INIT_56 => INIT_H_IDIG_56,
      INIT_57 => INIT_H_IDIG_57,
      INIT_58 => INIT_H_IDIG_58,
      INIT_59 => INIT_H_IDIG_59,
      INIT_5A => INIT_H_IDIG_5A,
      INIT_5B => INIT_H_IDIG_5B,
      INIT_5C => INIT_H_IDIG_5C,
      INIT_5D => INIT_H_IDIG_5D,
      INIT_5E => INIT_H_IDIG_5E,
      INIT_5F => INIT_H_IDIG_5F,
      INIT_60 => INIT_H_IDIG_60,
      INIT_61 => INIT_H_IDIG_61,
      INIT_62 => INIT_H_IDIG_62,
      INIT_63 => INIT_H_IDIG_63,
      INIT_64 => INIT_H_IDIG_64,
      INIT_65 => INIT_H_IDIG_65,
      INIT_66 => INIT_H_IDIG_66,
      INIT_67 => INIT_H_IDIG_67,
      INIT_68 => INIT_H_IDIG_68,
      INIT_69 => INIT_H_IDIG_69,
      INIT_6A => INIT_H_IDIG_6A,
      INIT_6B => INIT_H_IDIG_6B,
      INIT_6C => INIT_H_IDIG_6C,
      INIT_6D => INIT_H_IDIG_6D,
      INIT_6E => INIT_H_IDIG_6E,
      INIT_6F => INIT_H_IDIG_6F,
      INIT_70 => INIT_H_IDIG_70,
      INIT_71 => INIT_H_IDIG_71,
      INIT_72 => INIT_H_IDIG_72,
      INIT_73 => INIT_H_IDIG_73,
      INIT_74 => INIT_H_IDIG_74,
      INIT_75 => INIT_H_IDIG_75,
      INIT_76 => INIT_H_IDIG_76,
      INIT_77 => INIT_H_IDIG_77,
      INIT_78 => INIT_H_IDIG_78,
      INIT_79 => INIT_H_IDIG_79,
      INIT_7A => INIT_H_IDIG_7A,
      INIT_7B => INIT_H_IDIG_7B,
      INIT_7C => INIT_H_IDIG_7C,
      INIT_7D => INIT_H_IDIG_7D,
      INIT_7E => INIT_H_IDIG_7E,
      INIT_7F => INIT_H_IDIG_7F
   ) port map(
      ADDRARDADDR    => idig_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => idig_h_data_out_a(31 downto 0),
      DOPADOP        => idig_h_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );



   idig_l_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_L_IDIG_00,
      INIT_01 => INIT_L_IDIG_01,
      INIT_02 => INIT_L_IDIG_02,
      INIT_03 => INIT_L_IDIG_03,
      INIT_04 => INIT_L_IDIG_04,
      INIT_05 => INIT_L_IDIG_05,
      INIT_06 => INIT_L_IDIG_06,
      INIT_07 => INIT_L_IDIG_07,
      INIT_08 => INIT_L_IDIG_08,
      INIT_09 => INIT_L_IDIG_09,
      INIT_0A => INIT_L_IDIG_0A,
      INIT_0B => INIT_L_IDIG_0B,
      INIT_0C => INIT_L_IDIG_0C,
      INIT_0D => INIT_L_IDIG_0D,
      INIT_0E => INIT_L_IDIG_0E,
      INIT_0F => INIT_L_IDIG_0F,
      INIT_10 => INIT_L_IDIG_10,
      INIT_11 => INIT_L_IDIG_11,
      INIT_12 => INIT_L_IDIG_12,
      INIT_13 => INIT_L_IDIG_13,
      INIT_14 => INIT_L_IDIG_14,
      INIT_15 => INIT_L_IDIG_15,
      INIT_16 => INIT_L_IDIG_16,
      INIT_17 => INIT_L_IDIG_17,
      INIT_18 => INIT_L_IDIG_18,
      INIT_19 => INIT_L_IDIG_19,
      INIT_1A => INIT_L_IDIG_1A,
      INIT_1B => INIT_L_IDIG_1B,
      INIT_1C => INIT_L_IDIG_1C,
      INIT_1D => INIT_L_IDIG_1D,
      INIT_1E => INIT_L_IDIG_1E,
      INIT_1F => INIT_L_IDIG_1F,
      INIT_20 => INIT_L_IDIG_20,
      INIT_21 => INIT_L_IDIG_21,
      INIT_22 => INIT_L_IDIG_22,
      INIT_23 => INIT_L_IDIG_23,
      INIT_24 => INIT_L_IDIG_24,
      INIT_25 => INIT_L_IDIG_25,
      INIT_26 => INIT_L_IDIG_26,
      INIT_27 => INIT_L_IDIG_27,
      INIT_28 => INIT_L_IDIG_28,
      INIT_29 => INIT_L_IDIG_29,
      INIT_2A => INIT_L_IDIG_2A,
      INIT_2B => INIT_L_IDIG_2B,
      INIT_2C => INIT_L_IDIG_2C,
      INIT_2D => INIT_L_IDIG_2D,
      INIT_2E => INIT_L_IDIG_2E,
      INIT_2F => INIT_L_IDIG_2F,
      INIT_30 => INIT_L_IDIG_30,
      INIT_31 => INIT_L_IDIG_31,
      INIT_32 => INIT_L_IDIG_32,
      INIT_33 => INIT_L_IDIG_33,
      INIT_34 => INIT_L_IDIG_34,
      INIT_35 => INIT_L_IDIG_35,
      INIT_36 => INIT_L_IDIG_36,
      INIT_37 => INIT_L_IDIG_37,
      INIT_38 => INIT_L_IDIG_38,
      INIT_39 => INIT_L_IDIG_39,
      INIT_3A => INIT_L_IDIG_3A,
      INIT_3B => INIT_L_IDIG_3B,
      INIT_3C => INIT_L_IDIG_3C,
      INIT_3D => INIT_L_IDIG_3D,
      INIT_3E => INIT_L_IDIG_3E,
      INIT_3F => INIT_L_IDIG_3F,
      INIT_40 => INIT_L_IDIG_40,
      INIT_41 => INIT_L_IDIG_41,
      INIT_42 => INIT_L_IDIG_42,
      INIT_43 => INIT_L_IDIG_43,
      INIT_44 => INIT_L_IDIG_44,
      INIT_45 => INIT_L_IDIG_45,
      INIT_46 => INIT_L_IDIG_46,
      INIT_47 => INIT_L_IDIG_47,
      INIT_48 => INIT_L_IDIG_48,
      INIT_49 => INIT_L_IDIG_49,
      INIT_4A => INIT_L_IDIG_4A,
      INIT_4B => INIT_L_IDIG_4B,
      INIT_4C => INIT_L_IDIG_4C,
      INIT_4D => INIT_L_IDIG_4D,
      INIT_4E => INIT_L_IDIG_4E,
      INIT_4F => INIT_L_IDIG_4F,
      INIT_50 => INIT_L_IDIG_50,
      INIT_51 => INIT_L_IDIG_51,
      INIT_52 => INIT_L_IDIG_52,
      INIT_53 => INIT_L_IDIG_53,
      INIT_54 => INIT_L_IDIG_54,
      INIT_55 => INIT_L_IDIG_55,
      INIT_56 => INIT_L_IDIG_56,
      INIT_57 => INIT_L_IDIG_57,
      INIT_58 => INIT_L_IDIG_58,
      INIT_59 => INIT_L_IDIG_59,
      INIT_5A => INIT_L_IDIG_5A,
      INIT_5B => INIT_L_IDIG_5B,
      INIT_5C => INIT_L_IDIG_5C,
      INIT_5D => INIT_L_IDIG_5D,
      INIT_5E => INIT_L_IDIG_5E,
      INIT_5F => INIT_L_IDIG_5F,
      INIT_60 => INIT_L_IDIG_60,
      INIT_61 => INIT_L_IDIG_61,
      INIT_62 => INIT_L_IDIG_62,
      INIT_63 => INIT_L_IDIG_63,
      INIT_64 => INIT_L_IDIG_64,
      INIT_65 => INIT_L_IDIG_65,
      INIT_66 => INIT_L_IDIG_66,
      INIT_67 => INIT_L_IDIG_67,
      INIT_68 => INIT_L_IDIG_68,
      INIT_69 => INIT_L_IDIG_69,
      INIT_6A => INIT_L_IDIG_6A,
      INIT_6B => INIT_L_IDIG_6B,
      INIT_6C => INIT_L_IDIG_6C,
      INIT_6D => INIT_L_IDIG_6D,
      INIT_6E => INIT_L_IDIG_6E,
      INIT_6F => INIT_L_IDIG_6F,
      INIT_70 => INIT_L_IDIG_70,
      INIT_71 => INIT_L_IDIG_71,
      INIT_72 => INIT_L_IDIG_72,
      INIT_73 => INIT_L_IDIG_73,
      INIT_74 => INIT_L_IDIG_74,
      INIT_75 => INIT_L_IDIG_75,
      INIT_76 => INIT_L_IDIG_76,
      INIT_77 => INIT_L_IDIG_77,
      INIT_78 => INIT_L_IDIG_78,
      INIT_79 => INIT_L_IDIG_79,
      INIT_7A => INIT_L_IDIG_7A,
      INIT_7B => INIT_L_IDIG_7B,
      INIT_7C => INIT_L_IDIG_7C,
      INIT_7D => INIT_L_IDIG_7D,
      INIT_7E => INIT_L_IDIG_7E,
      INIT_7F => INIT_L_IDIG_7F
   ) port map(
      ADDRARDADDR    => idig_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => idig_l_data_out_a(31 downto 0),
      DOPADOP        => idig_l_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );

   idig_address_a <= '1' & adcData(4)(23 downto 12) & "111";
   outEnvData(4) <= x"0000" & idig_h_data_out_a(7 downto 0) & idig_l_data_out_a(7 downto 0);


   igua_h_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_H_IGUA_00,
      INIT_01 => INIT_H_IGUA_01,
      INIT_02 => INIT_H_IGUA_02,
      INIT_03 => INIT_H_IGUA_03,
      INIT_04 => INIT_H_IGUA_04,
      INIT_05 => INIT_H_IGUA_05,
      INIT_06 => INIT_H_IGUA_06,
      INIT_07 => INIT_H_IGUA_07,
      INIT_08 => INIT_H_IGUA_08,
      INIT_09 => INIT_H_IGUA_09,
      INIT_0A => INIT_H_IGUA_0A,
      INIT_0B => INIT_H_IGUA_0B,
      INIT_0C => INIT_H_IGUA_0C,
      INIT_0D => INIT_H_IGUA_0D,
      INIT_0E => INIT_H_IGUA_0E,
      INIT_0F => INIT_H_IGUA_0F,
      INIT_10 => INIT_H_IGUA_10,
      INIT_11 => INIT_H_IGUA_11,
      INIT_12 => INIT_H_IGUA_12,
      INIT_13 => INIT_H_IGUA_13,
      INIT_14 => INIT_H_IGUA_14,
      INIT_15 => INIT_H_IGUA_15,
      INIT_16 => INIT_H_IGUA_16,
      INIT_17 => INIT_H_IGUA_17,
      INIT_18 => INIT_H_IGUA_18,
      INIT_19 => INIT_H_IGUA_19,
      INIT_1A => INIT_H_IGUA_1A,
      INIT_1B => INIT_H_IGUA_1B,
      INIT_1C => INIT_H_IGUA_1C,
      INIT_1D => INIT_H_IGUA_1D,
      INIT_1E => INIT_H_IGUA_1E,
      INIT_1F => INIT_H_IGUA_1F,
      INIT_20 => INIT_H_IGUA_20,
      INIT_21 => INIT_H_IGUA_21,
      INIT_22 => INIT_H_IGUA_22,
      INIT_23 => INIT_H_IGUA_23,
      INIT_24 => INIT_H_IGUA_24,
      INIT_25 => INIT_H_IGUA_25,
      INIT_26 => INIT_H_IGUA_26,
      INIT_27 => INIT_H_IGUA_27,
      INIT_28 => INIT_H_IGUA_28,
      INIT_29 => INIT_H_IGUA_29,
      INIT_2A => INIT_H_IGUA_2A,
      INIT_2B => INIT_H_IGUA_2B,
      INIT_2C => INIT_H_IGUA_2C,
      INIT_2D => INIT_H_IGUA_2D,
      INIT_2E => INIT_H_IGUA_2E,
      INIT_2F => INIT_H_IGUA_2F,
      INIT_30 => INIT_H_IGUA_30,
      INIT_31 => INIT_H_IGUA_31,
      INIT_32 => INIT_H_IGUA_32,
      INIT_33 => INIT_H_IGUA_33,
      INIT_34 => INIT_H_IGUA_34,
      INIT_35 => INIT_H_IGUA_35,
      INIT_36 => INIT_H_IGUA_36,
      INIT_37 => INIT_H_IGUA_37,
      INIT_38 => INIT_H_IGUA_38,
      INIT_39 => INIT_H_IGUA_39,
      INIT_3A => INIT_H_IGUA_3A,
      INIT_3B => INIT_H_IGUA_3B,
      INIT_3C => INIT_H_IGUA_3C,
      INIT_3D => INIT_H_IGUA_3D,
      INIT_3E => INIT_H_IGUA_3E,
      INIT_3F => INIT_H_IGUA_3F,
      INIT_40 => INIT_H_IGUA_40,
      INIT_41 => INIT_H_IGUA_41,
      INIT_42 => INIT_H_IGUA_42,
      INIT_43 => INIT_H_IGUA_43,
      INIT_44 => INIT_H_IGUA_44,
      INIT_45 => INIT_H_IGUA_45,
      INIT_46 => INIT_H_IGUA_46,
      INIT_47 => INIT_H_IGUA_47,
      INIT_48 => INIT_H_IGUA_48,
      INIT_49 => INIT_H_IGUA_49,
      INIT_4A => INIT_H_IGUA_4A,
      INIT_4B => INIT_H_IGUA_4B,
      INIT_4C => INIT_H_IGUA_4C,
      INIT_4D => INIT_H_IGUA_4D,
      INIT_4E => INIT_H_IGUA_4E,
      INIT_4F => INIT_H_IGUA_4F,
      INIT_50 => INIT_H_IGUA_50,
      INIT_51 => INIT_H_IGUA_51,
      INIT_52 => INIT_H_IGUA_52,
      INIT_53 => INIT_H_IGUA_53,
      INIT_54 => INIT_H_IGUA_54,
      INIT_55 => INIT_H_IGUA_55,
      INIT_56 => INIT_H_IGUA_56,
      INIT_57 => INIT_H_IGUA_57,
      INIT_58 => INIT_H_IGUA_58,
      INIT_59 => INIT_H_IGUA_59,
      INIT_5A => INIT_H_IGUA_5A,
      INIT_5B => INIT_H_IGUA_5B,
      INIT_5C => INIT_H_IGUA_5C,
      INIT_5D => INIT_H_IGUA_5D,
      INIT_5E => INIT_H_IGUA_5E,
      INIT_5F => INIT_H_IGUA_5F,
      INIT_60 => INIT_H_IGUA_60,
      INIT_61 => INIT_H_IGUA_61,
      INIT_62 => INIT_H_IGUA_62,
      INIT_63 => INIT_H_IGUA_63,
      INIT_64 => INIT_H_IGUA_64,
      INIT_65 => INIT_H_IGUA_65,
      INIT_66 => INIT_H_IGUA_66,
      INIT_67 => INIT_H_IGUA_67,
      INIT_68 => INIT_H_IGUA_68,
      INIT_69 => INIT_H_IGUA_69,
      INIT_6A => INIT_H_IGUA_6A,
      INIT_6B => INIT_H_IGUA_6B,
      INIT_6C => INIT_H_IGUA_6C,
      INIT_6D => INIT_H_IGUA_6D,
      INIT_6E => INIT_H_IGUA_6E,
      INIT_6F => INIT_H_IGUA_6F,
      INIT_70 => INIT_H_IGUA_70,
      INIT_71 => INIT_H_IGUA_71,
      INIT_72 => INIT_H_IGUA_72,
      INIT_73 => INIT_H_IGUA_73,
      INIT_74 => INIT_H_IGUA_74,
      INIT_75 => INIT_H_IGUA_75,
      INIT_76 => INIT_H_IGUA_76,
      INIT_77 => INIT_H_IGUA_77,
      INIT_78 => INIT_H_IGUA_78,
      INIT_79 => INIT_H_IGUA_79,
      INIT_7A => INIT_H_IGUA_7A,
      INIT_7B => INIT_H_IGUA_7B,
      INIT_7C => INIT_H_IGUA_7C,
      INIT_7D => INIT_H_IGUA_7D,
      INIT_7E => INIT_H_IGUA_7E,
      INIT_7F => INIT_H_IGUA_7F
   ) port map(
      ADDRARDADDR    => igua_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => igua_h_data_out_a(31 downto 0),
      DOPADOP        => igua_h_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );



   igua_l_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_L_IGUA_00,
      INIT_01 => INIT_L_IGUA_01,
      INIT_02 => INIT_L_IGUA_02,
      INIT_03 => INIT_L_IGUA_03,
      INIT_04 => INIT_L_IGUA_04,
      INIT_05 => INIT_L_IGUA_05,
      INIT_06 => INIT_L_IGUA_06,
      INIT_07 => INIT_L_IGUA_07,
      INIT_08 => INIT_L_IGUA_08,
      INIT_09 => INIT_L_IGUA_09,
      INIT_0A => INIT_L_IGUA_0A,
      INIT_0B => INIT_L_IGUA_0B,
      INIT_0C => INIT_L_IGUA_0C,
      INIT_0D => INIT_L_IGUA_0D,
      INIT_0E => INIT_L_IGUA_0E,
      INIT_0F => INIT_L_IGUA_0F,
      INIT_10 => INIT_L_IGUA_10,
      INIT_11 => INIT_L_IGUA_11,
      INIT_12 => INIT_L_IGUA_12,
      INIT_13 => INIT_L_IGUA_13,
      INIT_14 => INIT_L_IGUA_14,
      INIT_15 => INIT_L_IGUA_15,
      INIT_16 => INIT_L_IGUA_16,
      INIT_17 => INIT_L_IGUA_17,
      INIT_18 => INIT_L_IGUA_18,
      INIT_19 => INIT_L_IGUA_19,
      INIT_1A => INIT_L_IGUA_1A,
      INIT_1B => INIT_L_IGUA_1B,
      INIT_1C => INIT_L_IGUA_1C,
      INIT_1D => INIT_L_IGUA_1D,
      INIT_1E => INIT_L_IGUA_1E,
      INIT_1F => INIT_L_IGUA_1F,
      INIT_20 => INIT_L_IGUA_20,
      INIT_21 => INIT_L_IGUA_21,
      INIT_22 => INIT_L_IGUA_22,
      INIT_23 => INIT_L_IGUA_23,
      INIT_24 => INIT_L_IGUA_24,
      INIT_25 => INIT_L_IGUA_25,
      INIT_26 => INIT_L_IGUA_26,
      INIT_27 => INIT_L_IGUA_27,
      INIT_28 => INIT_L_IGUA_28,
      INIT_29 => INIT_L_IGUA_29,
      INIT_2A => INIT_L_IGUA_2A,
      INIT_2B => INIT_L_IGUA_2B,
      INIT_2C => INIT_L_IGUA_2C,
      INIT_2D => INIT_L_IGUA_2D,
      INIT_2E => INIT_L_IGUA_2E,
      INIT_2F => INIT_L_IGUA_2F,
      INIT_30 => INIT_L_IGUA_30,
      INIT_31 => INIT_L_IGUA_31,
      INIT_32 => INIT_L_IGUA_32,
      INIT_33 => INIT_L_IGUA_33,
      INIT_34 => INIT_L_IGUA_34,
      INIT_35 => INIT_L_IGUA_35,
      INIT_36 => INIT_L_IGUA_36,
      INIT_37 => INIT_L_IGUA_37,
      INIT_38 => INIT_L_IGUA_38,
      INIT_39 => INIT_L_IGUA_39,
      INIT_3A => INIT_L_IGUA_3A,
      INIT_3B => INIT_L_IGUA_3B,
      INIT_3C => INIT_L_IGUA_3C,
      INIT_3D => INIT_L_IGUA_3D,
      INIT_3E => INIT_L_IGUA_3E,
      INIT_3F => INIT_L_IGUA_3F,
      INIT_40 => INIT_L_IGUA_40,
      INIT_41 => INIT_L_IGUA_41,
      INIT_42 => INIT_L_IGUA_42,
      INIT_43 => INIT_L_IGUA_43,
      INIT_44 => INIT_L_IGUA_44,
      INIT_45 => INIT_L_IGUA_45,
      INIT_46 => INIT_L_IGUA_46,
      INIT_47 => INIT_L_IGUA_47,
      INIT_48 => INIT_L_IGUA_48,
      INIT_49 => INIT_L_IGUA_49,
      INIT_4A => INIT_L_IGUA_4A,
      INIT_4B => INIT_L_IGUA_4B,
      INIT_4C => INIT_L_IGUA_4C,
      INIT_4D => INIT_L_IGUA_4D,
      INIT_4E => INIT_L_IGUA_4E,
      INIT_4F => INIT_L_IGUA_4F,
      INIT_50 => INIT_L_IGUA_50,
      INIT_51 => INIT_L_IGUA_51,
      INIT_52 => INIT_L_IGUA_52,
      INIT_53 => INIT_L_IGUA_53,
      INIT_54 => INIT_L_IGUA_54,
      INIT_55 => INIT_L_IGUA_55,
      INIT_56 => INIT_L_IGUA_56,
      INIT_57 => INIT_L_IGUA_57,
      INIT_58 => INIT_L_IGUA_58,
      INIT_59 => INIT_L_IGUA_59,
      INIT_5A => INIT_L_IGUA_5A,
      INIT_5B => INIT_L_IGUA_5B,
      INIT_5C => INIT_L_IGUA_5C,
      INIT_5D => INIT_L_IGUA_5D,
      INIT_5E => INIT_L_IGUA_5E,
      INIT_5F => INIT_L_IGUA_5F,
      INIT_60 => INIT_L_IGUA_60,
      INIT_61 => INIT_L_IGUA_61,
      INIT_62 => INIT_L_IGUA_62,
      INIT_63 => INIT_L_IGUA_63,
      INIT_64 => INIT_L_IGUA_64,
      INIT_65 => INIT_L_IGUA_65,
      INIT_66 => INIT_L_IGUA_66,
      INIT_67 => INIT_L_IGUA_67,
      INIT_68 => INIT_L_IGUA_68,
      INIT_69 => INIT_L_IGUA_69,
      INIT_6A => INIT_L_IGUA_6A,
      INIT_6B => INIT_L_IGUA_6B,
      INIT_6C => INIT_L_IGUA_6C,
      INIT_6D => INIT_L_IGUA_6D,
      INIT_6E => INIT_L_IGUA_6E,
      INIT_6F => INIT_L_IGUA_6F,
      INIT_70 => INIT_L_IGUA_70,
      INIT_71 => INIT_L_IGUA_71,
      INIT_72 => INIT_L_IGUA_72,
      INIT_73 => INIT_L_IGUA_73,
      INIT_74 => INIT_L_IGUA_74,
      INIT_75 => INIT_L_IGUA_75,
      INIT_76 => INIT_L_IGUA_76,
      INIT_77 => INIT_L_IGUA_77,
      INIT_78 => INIT_L_IGUA_78,
      INIT_79 => INIT_L_IGUA_79,
      INIT_7A => INIT_L_IGUA_7A,
      INIT_7B => INIT_L_IGUA_7B,
      INIT_7C => INIT_L_IGUA_7C,
      INIT_7D => INIT_L_IGUA_7D,
      INIT_7E => INIT_L_IGUA_7E,
      INIT_7F => INIT_L_IGUA_7F
   ) port map(
      ADDRARDADDR    => igua_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => igua_l_data_out_a(31 downto 0),
      DOPADOP        => igua_l_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );

   igua_address_a <= '1' & adcData(5)(23 downto 12) & "111";
   outEnvData(5) <= x"0000" & igua_h_data_out_a(7 downto 0) & igua_l_data_out_a(7 downto 0);


   ibia_h_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_H_IBIA_00,
      INIT_01 => INIT_H_IBIA_01,
      INIT_02 => INIT_H_IBIA_02,
      INIT_03 => INIT_H_IBIA_03,
      INIT_04 => INIT_H_IBIA_04,
      INIT_05 => INIT_H_IBIA_05,
      INIT_06 => INIT_H_IBIA_06,
      INIT_07 => INIT_H_IBIA_07,
      INIT_08 => INIT_H_IBIA_08,
      INIT_09 => INIT_H_IBIA_09,
      INIT_0A => INIT_H_IBIA_0A,
      INIT_0B => INIT_H_IBIA_0B,
      INIT_0C => INIT_H_IBIA_0C,
      INIT_0D => INIT_H_IBIA_0D,
      INIT_0E => INIT_H_IBIA_0E,
      INIT_0F => INIT_H_IBIA_0F,
      INIT_10 => INIT_H_IBIA_10,
      INIT_11 => INIT_H_IBIA_11,
      INIT_12 => INIT_H_IBIA_12,
      INIT_13 => INIT_H_IBIA_13,
      INIT_14 => INIT_H_IBIA_14,
      INIT_15 => INIT_H_IBIA_15,
      INIT_16 => INIT_H_IBIA_16,
      INIT_17 => INIT_H_IBIA_17,
      INIT_18 => INIT_H_IBIA_18,
      INIT_19 => INIT_H_IBIA_19,
      INIT_1A => INIT_H_IBIA_1A,
      INIT_1B => INIT_H_IBIA_1B,
      INIT_1C => INIT_H_IBIA_1C,
      INIT_1D => INIT_H_IBIA_1D,
      INIT_1E => INIT_H_IBIA_1E,
      INIT_1F => INIT_H_IBIA_1F,
      INIT_20 => INIT_H_IBIA_20,
      INIT_21 => INIT_H_IBIA_21,
      INIT_22 => INIT_H_IBIA_22,
      INIT_23 => INIT_H_IBIA_23,
      INIT_24 => INIT_H_IBIA_24,
      INIT_25 => INIT_H_IBIA_25,
      INIT_26 => INIT_H_IBIA_26,
      INIT_27 => INIT_H_IBIA_27,
      INIT_28 => INIT_H_IBIA_28,
      INIT_29 => INIT_H_IBIA_29,
      INIT_2A => INIT_H_IBIA_2A,
      INIT_2B => INIT_H_IBIA_2B,
      INIT_2C => INIT_H_IBIA_2C,
      INIT_2D => INIT_H_IBIA_2D,
      INIT_2E => INIT_H_IBIA_2E,
      INIT_2F => INIT_H_IBIA_2F,
      INIT_30 => INIT_H_IBIA_30,
      INIT_31 => INIT_H_IBIA_31,
      INIT_32 => INIT_H_IBIA_32,
      INIT_33 => INIT_H_IBIA_33,
      INIT_34 => INIT_H_IBIA_34,
      INIT_35 => INIT_H_IBIA_35,
      INIT_36 => INIT_H_IBIA_36,
      INIT_37 => INIT_H_IBIA_37,
      INIT_38 => INIT_H_IBIA_38,
      INIT_39 => INIT_H_IBIA_39,
      INIT_3A => INIT_H_IBIA_3A,
      INIT_3B => INIT_H_IBIA_3B,
      INIT_3C => INIT_H_IBIA_3C,
      INIT_3D => INIT_H_IBIA_3D,
      INIT_3E => INIT_H_IBIA_3E,
      INIT_3F => INIT_H_IBIA_3F,
      INIT_40 => INIT_H_IBIA_40,
      INIT_41 => INIT_H_IBIA_41,
      INIT_42 => INIT_H_IBIA_42,
      INIT_43 => INIT_H_IBIA_43,
      INIT_44 => INIT_H_IBIA_44,
      INIT_45 => INIT_H_IBIA_45,
      INIT_46 => INIT_H_IBIA_46,
      INIT_47 => INIT_H_IBIA_47,
      INIT_48 => INIT_H_IBIA_48,
      INIT_49 => INIT_H_IBIA_49,
      INIT_4A => INIT_H_IBIA_4A,
      INIT_4B => INIT_H_IBIA_4B,
      INIT_4C => INIT_H_IBIA_4C,
      INIT_4D => INIT_H_IBIA_4D,
      INIT_4E => INIT_H_IBIA_4E,
      INIT_4F => INIT_H_IBIA_4F,
      INIT_50 => INIT_H_IBIA_50,
      INIT_51 => INIT_H_IBIA_51,
      INIT_52 => INIT_H_IBIA_52,
      INIT_53 => INIT_H_IBIA_53,
      INIT_54 => INIT_H_IBIA_54,
      INIT_55 => INIT_H_IBIA_55,
      INIT_56 => INIT_H_IBIA_56,
      INIT_57 => INIT_H_IBIA_57,
      INIT_58 => INIT_H_IBIA_58,
      INIT_59 => INIT_H_IBIA_59,
      INIT_5A => INIT_H_IBIA_5A,
      INIT_5B => INIT_H_IBIA_5B,
      INIT_5C => INIT_H_IBIA_5C,
      INIT_5D => INIT_H_IBIA_5D,
      INIT_5E => INIT_H_IBIA_5E,
      INIT_5F => INIT_H_IBIA_5F,
      INIT_60 => INIT_H_IBIA_60,
      INIT_61 => INIT_H_IBIA_61,
      INIT_62 => INIT_H_IBIA_62,
      INIT_63 => INIT_H_IBIA_63,
      INIT_64 => INIT_H_IBIA_64,
      INIT_65 => INIT_H_IBIA_65,
      INIT_66 => INIT_H_IBIA_66,
      INIT_67 => INIT_H_IBIA_67,
      INIT_68 => INIT_H_IBIA_68,
      INIT_69 => INIT_H_IBIA_69,
      INIT_6A => INIT_H_IBIA_6A,
      INIT_6B => INIT_H_IBIA_6B,
      INIT_6C => INIT_H_IBIA_6C,
      INIT_6D => INIT_H_IBIA_6D,
      INIT_6E => INIT_H_IBIA_6E,
      INIT_6F => INIT_H_IBIA_6F,
      INIT_70 => INIT_H_IBIA_70,
      INIT_71 => INIT_H_IBIA_71,
      INIT_72 => INIT_H_IBIA_72,
      INIT_73 => INIT_H_IBIA_73,
      INIT_74 => INIT_H_IBIA_74,
      INIT_75 => INIT_H_IBIA_75,
      INIT_76 => INIT_H_IBIA_76,
      INIT_77 => INIT_H_IBIA_77,
      INIT_78 => INIT_H_IBIA_78,
      INIT_79 => INIT_H_IBIA_79,
      INIT_7A => INIT_H_IBIA_7A,
      INIT_7B => INIT_H_IBIA_7B,
      INIT_7C => INIT_H_IBIA_7C,
      INIT_7D => INIT_H_IBIA_7D,
      INIT_7E => INIT_H_IBIA_7E,
      INIT_7F => INIT_H_IBIA_7F
   ) port map(
      ADDRARDADDR    => ibia_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => ibia_h_data_out_a(31 downto 0),
      DOPADOP        => ibia_h_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );



   ibia_l_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_L_IBIA_00,
      INIT_01 => INIT_L_IBIA_01,
      INIT_02 => INIT_L_IBIA_02,
      INIT_03 => INIT_L_IBIA_03,
      INIT_04 => INIT_L_IBIA_04,
      INIT_05 => INIT_L_IBIA_05,
      INIT_06 => INIT_L_IBIA_06,
      INIT_07 => INIT_L_IBIA_07,
      INIT_08 => INIT_L_IBIA_08,
      INIT_09 => INIT_L_IBIA_09,
      INIT_0A => INIT_L_IBIA_0A,
      INIT_0B => INIT_L_IBIA_0B,
      INIT_0C => INIT_L_IBIA_0C,
      INIT_0D => INIT_L_IBIA_0D,
      INIT_0E => INIT_L_IBIA_0E,
      INIT_0F => INIT_L_IBIA_0F,
      INIT_10 => INIT_L_IBIA_10,
      INIT_11 => INIT_L_IBIA_11,
      INIT_12 => INIT_L_IBIA_12,
      INIT_13 => INIT_L_IBIA_13,
      INIT_14 => INIT_L_IBIA_14,
      INIT_15 => INIT_L_IBIA_15,
      INIT_16 => INIT_L_IBIA_16,
      INIT_17 => INIT_L_IBIA_17,
      INIT_18 => INIT_L_IBIA_18,
      INIT_19 => INIT_L_IBIA_19,
      INIT_1A => INIT_L_IBIA_1A,
      INIT_1B => INIT_L_IBIA_1B,
      INIT_1C => INIT_L_IBIA_1C,
      INIT_1D => INIT_L_IBIA_1D,
      INIT_1E => INIT_L_IBIA_1E,
      INIT_1F => INIT_L_IBIA_1F,
      INIT_20 => INIT_L_IBIA_20,
      INIT_21 => INIT_L_IBIA_21,
      INIT_22 => INIT_L_IBIA_22,
      INIT_23 => INIT_L_IBIA_23,
      INIT_24 => INIT_L_IBIA_24,
      INIT_25 => INIT_L_IBIA_25,
      INIT_26 => INIT_L_IBIA_26,
      INIT_27 => INIT_L_IBIA_27,
      INIT_28 => INIT_L_IBIA_28,
      INIT_29 => INIT_L_IBIA_29,
      INIT_2A => INIT_L_IBIA_2A,
      INIT_2B => INIT_L_IBIA_2B,
      INIT_2C => INIT_L_IBIA_2C,
      INIT_2D => INIT_L_IBIA_2D,
      INIT_2E => INIT_L_IBIA_2E,
      INIT_2F => INIT_L_IBIA_2F,
      INIT_30 => INIT_L_IBIA_30,
      INIT_31 => INIT_L_IBIA_31,
      INIT_32 => INIT_L_IBIA_32,
      INIT_33 => INIT_L_IBIA_33,
      INIT_34 => INIT_L_IBIA_34,
      INIT_35 => INIT_L_IBIA_35,
      INIT_36 => INIT_L_IBIA_36,
      INIT_37 => INIT_L_IBIA_37,
      INIT_38 => INIT_L_IBIA_38,
      INIT_39 => INIT_L_IBIA_39,
      INIT_3A => INIT_L_IBIA_3A,
      INIT_3B => INIT_L_IBIA_3B,
      INIT_3C => INIT_L_IBIA_3C,
      INIT_3D => INIT_L_IBIA_3D,
      INIT_3E => INIT_L_IBIA_3E,
      INIT_3F => INIT_L_IBIA_3F,
      INIT_40 => INIT_L_IBIA_40,
      INIT_41 => INIT_L_IBIA_41,
      INIT_42 => INIT_L_IBIA_42,
      INIT_43 => INIT_L_IBIA_43,
      INIT_44 => INIT_L_IBIA_44,
      INIT_45 => INIT_L_IBIA_45,
      INIT_46 => INIT_L_IBIA_46,
      INIT_47 => INIT_L_IBIA_47,
      INIT_48 => INIT_L_IBIA_48,
      INIT_49 => INIT_L_IBIA_49,
      INIT_4A => INIT_L_IBIA_4A,
      INIT_4B => INIT_L_IBIA_4B,
      INIT_4C => INIT_L_IBIA_4C,
      INIT_4D => INIT_L_IBIA_4D,
      INIT_4E => INIT_L_IBIA_4E,
      INIT_4F => INIT_L_IBIA_4F,
      INIT_50 => INIT_L_IBIA_50,
      INIT_51 => INIT_L_IBIA_51,
      INIT_52 => INIT_L_IBIA_52,
      INIT_53 => INIT_L_IBIA_53,
      INIT_54 => INIT_L_IBIA_54,
      INIT_55 => INIT_L_IBIA_55,
      INIT_56 => INIT_L_IBIA_56,
      INIT_57 => INIT_L_IBIA_57,
      INIT_58 => INIT_L_IBIA_58,
      INIT_59 => INIT_L_IBIA_59,
      INIT_5A => INIT_L_IBIA_5A,
      INIT_5B => INIT_L_IBIA_5B,
      INIT_5C => INIT_L_IBIA_5C,
      INIT_5D => INIT_L_IBIA_5D,
      INIT_5E => INIT_L_IBIA_5E,
      INIT_5F => INIT_L_IBIA_5F,
      INIT_60 => INIT_L_IBIA_60,
      INIT_61 => INIT_L_IBIA_61,
      INIT_62 => INIT_L_IBIA_62,
      INIT_63 => INIT_L_IBIA_63,
      INIT_64 => INIT_L_IBIA_64,
      INIT_65 => INIT_L_IBIA_65,
      INIT_66 => INIT_L_IBIA_66,
      INIT_67 => INIT_L_IBIA_67,
      INIT_68 => INIT_L_IBIA_68,
      INIT_69 => INIT_L_IBIA_69,
      INIT_6A => INIT_L_IBIA_6A,
      INIT_6B => INIT_L_IBIA_6B,
      INIT_6C => INIT_L_IBIA_6C,
      INIT_6D => INIT_L_IBIA_6D,
      INIT_6E => INIT_L_IBIA_6E,
      INIT_6F => INIT_L_IBIA_6F,
      INIT_70 => INIT_L_IBIA_70,
      INIT_71 => INIT_L_IBIA_71,
      INIT_72 => INIT_L_IBIA_72,
      INIT_73 => INIT_L_IBIA_73,
      INIT_74 => INIT_L_IBIA_74,
      INIT_75 => INIT_L_IBIA_75,
      INIT_76 => INIT_L_IBIA_76,
      INIT_77 => INIT_L_IBIA_77,
      INIT_78 => INIT_L_IBIA_78,
      INIT_79 => INIT_L_IBIA_79,
      INIT_7A => INIT_L_IBIA_7A,
      INIT_7B => INIT_L_IBIA_7B,
      INIT_7C => INIT_L_IBIA_7C,
      INIT_7D => INIT_L_IBIA_7D,
      INIT_7E => INIT_L_IBIA_7E,
      INIT_7F => INIT_L_IBIA_7F
   ) port map(
      ADDRARDADDR    => ibia_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => ibia_l_data_out_a(31 downto 0),
      DOPADOP        => ibia_l_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );

   ibia_address_a <= '1' & adcData(6)(23 downto 12) & "111";
   outEnvData(6) <= x"0000" & ibia_h_data_out_a(7 downto 0) & ibia_l_data_out_a(7 downto 0);


   avin_h_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_H_AVIN_00,
      INIT_01 => INIT_H_AVIN_01,
      INIT_02 => INIT_H_AVIN_02,
      INIT_03 => INIT_H_AVIN_03,
      INIT_04 => INIT_H_AVIN_04,
      INIT_05 => INIT_H_AVIN_05,
      INIT_06 => INIT_H_AVIN_06,
      INIT_07 => INIT_H_AVIN_07,
      INIT_08 => INIT_H_AVIN_08,
      INIT_09 => INIT_H_AVIN_09,
      INIT_0A => INIT_H_AVIN_0A,
      INIT_0B => INIT_H_AVIN_0B,
      INIT_0C => INIT_H_AVIN_0C,
      INIT_0D => INIT_H_AVIN_0D,
      INIT_0E => INIT_H_AVIN_0E,
      INIT_0F => INIT_H_AVIN_0F,
      INIT_10 => INIT_H_AVIN_10,
      INIT_11 => INIT_H_AVIN_11,
      INIT_12 => INIT_H_AVIN_12,
      INIT_13 => INIT_H_AVIN_13,
      INIT_14 => INIT_H_AVIN_14,
      INIT_15 => INIT_H_AVIN_15,
      INIT_16 => INIT_H_AVIN_16,
      INIT_17 => INIT_H_AVIN_17,
      INIT_18 => INIT_H_AVIN_18,
      INIT_19 => INIT_H_AVIN_19,
      INIT_1A => INIT_H_AVIN_1A,
      INIT_1B => INIT_H_AVIN_1B,
      INIT_1C => INIT_H_AVIN_1C,
      INIT_1D => INIT_H_AVIN_1D,
      INIT_1E => INIT_H_AVIN_1E,
      INIT_1F => INIT_H_AVIN_1F,
      INIT_20 => INIT_H_AVIN_20,
      INIT_21 => INIT_H_AVIN_21,
      INIT_22 => INIT_H_AVIN_22,
      INIT_23 => INIT_H_AVIN_23,
      INIT_24 => INIT_H_AVIN_24,
      INIT_25 => INIT_H_AVIN_25,
      INIT_26 => INIT_H_AVIN_26,
      INIT_27 => INIT_H_AVIN_27,
      INIT_28 => INIT_H_AVIN_28,
      INIT_29 => INIT_H_AVIN_29,
      INIT_2A => INIT_H_AVIN_2A,
      INIT_2B => INIT_H_AVIN_2B,
      INIT_2C => INIT_H_AVIN_2C,
      INIT_2D => INIT_H_AVIN_2D,
      INIT_2E => INIT_H_AVIN_2E,
      INIT_2F => INIT_H_AVIN_2F,
      INIT_30 => INIT_H_AVIN_30,
      INIT_31 => INIT_H_AVIN_31,
      INIT_32 => INIT_H_AVIN_32,
      INIT_33 => INIT_H_AVIN_33,
      INIT_34 => INIT_H_AVIN_34,
      INIT_35 => INIT_H_AVIN_35,
      INIT_36 => INIT_H_AVIN_36,
      INIT_37 => INIT_H_AVIN_37,
      INIT_38 => INIT_H_AVIN_38,
      INIT_39 => INIT_H_AVIN_39,
      INIT_3A => INIT_H_AVIN_3A,
      INIT_3B => INIT_H_AVIN_3B,
      INIT_3C => INIT_H_AVIN_3C,
      INIT_3D => INIT_H_AVIN_3D,
      INIT_3E => INIT_H_AVIN_3E,
      INIT_3F => INIT_H_AVIN_3F,
      INIT_40 => INIT_H_AVIN_40,
      INIT_41 => INIT_H_AVIN_41,
      INIT_42 => INIT_H_AVIN_42,
      INIT_43 => INIT_H_AVIN_43,
      INIT_44 => INIT_H_AVIN_44,
      INIT_45 => INIT_H_AVIN_45,
      INIT_46 => INIT_H_AVIN_46,
      INIT_47 => INIT_H_AVIN_47,
      INIT_48 => INIT_H_AVIN_48,
      INIT_49 => INIT_H_AVIN_49,
      INIT_4A => INIT_H_AVIN_4A,
      INIT_4B => INIT_H_AVIN_4B,
      INIT_4C => INIT_H_AVIN_4C,
      INIT_4D => INIT_H_AVIN_4D,
      INIT_4E => INIT_H_AVIN_4E,
      INIT_4F => INIT_H_AVIN_4F,
      INIT_50 => INIT_H_AVIN_50,
      INIT_51 => INIT_H_AVIN_51,
      INIT_52 => INIT_H_AVIN_52,
      INIT_53 => INIT_H_AVIN_53,
      INIT_54 => INIT_H_AVIN_54,
      INIT_55 => INIT_H_AVIN_55,
      INIT_56 => INIT_H_AVIN_56,
      INIT_57 => INIT_H_AVIN_57,
      INIT_58 => INIT_H_AVIN_58,
      INIT_59 => INIT_H_AVIN_59,
      INIT_5A => INIT_H_AVIN_5A,
      INIT_5B => INIT_H_AVIN_5B,
      INIT_5C => INIT_H_AVIN_5C,
      INIT_5D => INIT_H_AVIN_5D,
      INIT_5E => INIT_H_AVIN_5E,
      INIT_5F => INIT_H_AVIN_5F,
      INIT_60 => INIT_H_AVIN_60,
      INIT_61 => INIT_H_AVIN_61,
      INIT_62 => INIT_H_AVIN_62,
      INIT_63 => INIT_H_AVIN_63,
      INIT_64 => INIT_H_AVIN_64,
      INIT_65 => INIT_H_AVIN_65,
      INIT_66 => INIT_H_AVIN_66,
      INIT_67 => INIT_H_AVIN_67,
      INIT_68 => INIT_H_AVIN_68,
      INIT_69 => INIT_H_AVIN_69,
      INIT_6A => INIT_H_AVIN_6A,
      INIT_6B => INIT_H_AVIN_6B,
      INIT_6C => INIT_H_AVIN_6C,
      INIT_6D => INIT_H_AVIN_6D,
      INIT_6E => INIT_H_AVIN_6E,
      INIT_6F => INIT_H_AVIN_6F,
      INIT_70 => INIT_H_AVIN_70,
      INIT_71 => INIT_H_AVIN_71,
      INIT_72 => INIT_H_AVIN_72,
      INIT_73 => INIT_H_AVIN_73,
      INIT_74 => INIT_H_AVIN_74,
      INIT_75 => INIT_H_AVIN_75,
      INIT_76 => INIT_H_AVIN_76,
      INIT_77 => INIT_H_AVIN_77,
      INIT_78 => INIT_H_AVIN_78,
      INIT_79 => INIT_H_AVIN_79,
      INIT_7A => INIT_H_AVIN_7A,
      INIT_7B => INIT_H_AVIN_7B,
      INIT_7C => INIT_H_AVIN_7C,
      INIT_7D => INIT_H_AVIN_7D,
      INIT_7E => INIT_H_AVIN_7E,
      INIT_7F => INIT_H_AVIN_7F
   ) port map(
      ADDRARDADDR    => avin_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => avin_h_data_out_a(31 downto 0),
      DOPADOP        => avin_h_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );



   avin_l_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_L_AVIN_00,
      INIT_01 => INIT_L_AVIN_01,
      INIT_02 => INIT_L_AVIN_02,
      INIT_03 => INIT_L_AVIN_03,
      INIT_04 => INIT_L_AVIN_04,
      INIT_05 => INIT_L_AVIN_05,
      INIT_06 => INIT_L_AVIN_06,
      INIT_07 => INIT_L_AVIN_07,
      INIT_08 => INIT_L_AVIN_08,
      INIT_09 => INIT_L_AVIN_09,
      INIT_0A => INIT_L_AVIN_0A,
      INIT_0B => INIT_L_AVIN_0B,
      INIT_0C => INIT_L_AVIN_0C,
      INIT_0D => INIT_L_AVIN_0D,
      INIT_0E => INIT_L_AVIN_0E,
      INIT_0F => INIT_L_AVIN_0F,
      INIT_10 => INIT_L_AVIN_10,
      INIT_11 => INIT_L_AVIN_11,
      INIT_12 => INIT_L_AVIN_12,
      INIT_13 => INIT_L_AVIN_13,
      INIT_14 => INIT_L_AVIN_14,
      INIT_15 => INIT_L_AVIN_15,
      INIT_16 => INIT_L_AVIN_16,
      INIT_17 => INIT_L_AVIN_17,
      INIT_18 => INIT_L_AVIN_18,
      INIT_19 => INIT_L_AVIN_19,
      INIT_1A => INIT_L_AVIN_1A,
      INIT_1B => INIT_L_AVIN_1B,
      INIT_1C => INIT_L_AVIN_1C,
      INIT_1D => INIT_L_AVIN_1D,
      INIT_1E => INIT_L_AVIN_1E,
      INIT_1F => INIT_L_AVIN_1F,
      INIT_20 => INIT_L_AVIN_20,
      INIT_21 => INIT_L_AVIN_21,
      INIT_22 => INIT_L_AVIN_22,
      INIT_23 => INIT_L_AVIN_23,
      INIT_24 => INIT_L_AVIN_24,
      INIT_25 => INIT_L_AVIN_25,
      INIT_26 => INIT_L_AVIN_26,
      INIT_27 => INIT_L_AVIN_27,
      INIT_28 => INIT_L_AVIN_28,
      INIT_29 => INIT_L_AVIN_29,
      INIT_2A => INIT_L_AVIN_2A,
      INIT_2B => INIT_L_AVIN_2B,
      INIT_2C => INIT_L_AVIN_2C,
      INIT_2D => INIT_L_AVIN_2D,
      INIT_2E => INIT_L_AVIN_2E,
      INIT_2F => INIT_L_AVIN_2F,
      INIT_30 => INIT_L_AVIN_30,
      INIT_31 => INIT_L_AVIN_31,
      INIT_32 => INIT_L_AVIN_32,
      INIT_33 => INIT_L_AVIN_33,
      INIT_34 => INIT_L_AVIN_34,
      INIT_35 => INIT_L_AVIN_35,
      INIT_36 => INIT_L_AVIN_36,
      INIT_37 => INIT_L_AVIN_37,
      INIT_38 => INIT_L_AVIN_38,
      INIT_39 => INIT_L_AVIN_39,
      INIT_3A => INIT_L_AVIN_3A,
      INIT_3B => INIT_L_AVIN_3B,
      INIT_3C => INIT_L_AVIN_3C,
      INIT_3D => INIT_L_AVIN_3D,
      INIT_3E => INIT_L_AVIN_3E,
      INIT_3F => INIT_L_AVIN_3F,
      INIT_40 => INIT_L_AVIN_40,
      INIT_41 => INIT_L_AVIN_41,
      INIT_42 => INIT_L_AVIN_42,
      INIT_43 => INIT_L_AVIN_43,
      INIT_44 => INIT_L_AVIN_44,
      INIT_45 => INIT_L_AVIN_45,
      INIT_46 => INIT_L_AVIN_46,
      INIT_47 => INIT_L_AVIN_47,
      INIT_48 => INIT_L_AVIN_48,
      INIT_49 => INIT_L_AVIN_49,
      INIT_4A => INIT_L_AVIN_4A,
      INIT_4B => INIT_L_AVIN_4B,
      INIT_4C => INIT_L_AVIN_4C,
      INIT_4D => INIT_L_AVIN_4D,
      INIT_4E => INIT_L_AVIN_4E,
      INIT_4F => INIT_L_AVIN_4F,
      INIT_50 => INIT_L_AVIN_50,
      INIT_51 => INIT_L_AVIN_51,
      INIT_52 => INIT_L_AVIN_52,
      INIT_53 => INIT_L_AVIN_53,
      INIT_54 => INIT_L_AVIN_54,
      INIT_55 => INIT_L_AVIN_55,
      INIT_56 => INIT_L_AVIN_56,
      INIT_57 => INIT_L_AVIN_57,
      INIT_58 => INIT_L_AVIN_58,
      INIT_59 => INIT_L_AVIN_59,
      INIT_5A => INIT_L_AVIN_5A,
      INIT_5B => INIT_L_AVIN_5B,
      INIT_5C => INIT_L_AVIN_5C,
      INIT_5D => INIT_L_AVIN_5D,
      INIT_5E => INIT_L_AVIN_5E,
      INIT_5F => INIT_L_AVIN_5F,
      INIT_60 => INIT_L_AVIN_60,
      INIT_61 => INIT_L_AVIN_61,
      INIT_62 => INIT_L_AVIN_62,
      INIT_63 => INIT_L_AVIN_63,
      INIT_64 => INIT_L_AVIN_64,
      INIT_65 => INIT_L_AVIN_65,
      INIT_66 => INIT_L_AVIN_66,
      INIT_67 => INIT_L_AVIN_67,
      INIT_68 => INIT_L_AVIN_68,
      INIT_69 => INIT_L_AVIN_69,
      INIT_6A => INIT_L_AVIN_6A,
      INIT_6B => INIT_L_AVIN_6B,
      INIT_6C => INIT_L_AVIN_6C,
      INIT_6D => INIT_L_AVIN_6D,
      INIT_6E => INIT_L_AVIN_6E,
      INIT_6F => INIT_L_AVIN_6F,
      INIT_70 => INIT_L_AVIN_70,
      INIT_71 => INIT_L_AVIN_71,
      INIT_72 => INIT_L_AVIN_72,
      INIT_73 => INIT_L_AVIN_73,
      INIT_74 => INIT_L_AVIN_74,
      INIT_75 => INIT_L_AVIN_75,
      INIT_76 => INIT_L_AVIN_76,
      INIT_77 => INIT_L_AVIN_77,
      INIT_78 => INIT_L_AVIN_78,
      INIT_79 => INIT_L_AVIN_79,
      INIT_7A => INIT_L_AVIN_7A,
      INIT_7B => INIT_L_AVIN_7B,
      INIT_7C => INIT_L_AVIN_7C,
      INIT_7D => INIT_L_AVIN_7D,
      INIT_7E => INIT_L_AVIN_7E,
      INIT_7F => INIT_L_AVIN_7F
   ) port map(
      ADDRARDADDR    => avin_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => avin_l_data_out_a(31 downto 0),
      DOPADOP        => avin_l_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );

   avin_address_a <= '1' & adcData(7)(23 downto 12) & "111";
   outEnvData(7) <= x"0000" & avin_h_data_out_a(7 downto 0) & avin_l_data_out_a(7 downto 0);


   dvin_h_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_H_DVIN_00,
      INIT_01 => INIT_H_DVIN_01,
      INIT_02 => INIT_H_DVIN_02,
      INIT_03 => INIT_H_DVIN_03,
      INIT_04 => INIT_H_DVIN_04,
      INIT_05 => INIT_H_DVIN_05,
      INIT_06 => INIT_H_DVIN_06,
      INIT_07 => INIT_H_DVIN_07,
      INIT_08 => INIT_H_DVIN_08,
      INIT_09 => INIT_H_DVIN_09,
      INIT_0A => INIT_H_DVIN_0A,
      INIT_0B => INIT_H_DVIN_0B,
      INIT_0C => INIT_H_DVIN_0C,
      INIT_0D => INIT_H_DVIN_0D,
      INIT_0E => INIT_H_DVIN_0E,
      INIT_0F => INIT_H_DVIN_0F,
      INIT_10 => INIT_H_DVIN_10,
      INIT_11 => INIT_H_DVIN_11,
      INIT_12 => INIT_H_DVIN_12,
      INIT_13 => INIT_H_DVIN_13,
      INIT_14 => INIT_H_DVIN_14,
      INIT_15 => INIT_H_DVIN_15,
      INIT_16 => INIT_H_DVIN_16,
      INIT_17 => INIT_H_DVIN_17,
      INIT_18 => INIT_H_DVIN_18,
      INIT_19 => INIT_H_DVIN_19,
      INIT_1A => INIT_H_DVIN_1A,
      INIT_1B => INIT_H_DVIN_1B,
      INIT_1C => INIT_H_DVIN_1C,
      INIT_1D => INIT_H_DVIN_1D,
      INIT_1E => INIT_H_DVIN_1E,
      INIT_1F => INIT_H_DVIN_1F,
      INIT_20 => INIT_H_DVIN_20,
      INIT_21 => INIT_H_DVIN_21,
      INIT_22 => INIT_H_DVIN_22,
      INIT_23 => INIT_H_DVIN_23,
      INIT_24 => INIT_H_DVIN_24,
      INIT_25 => INIT_H_DVIN_25,
      INIT_26 => INIT_H_DVIN_26,
      INIT_27 => INIT_H_DVIN_27,
      INIT_28 => INIT_H_DVIN_28,
      INIT_29 => INIT_H_DVIN_29,
      INIT_2A => INIT_H_DVIN_2A,
      INIT_2B => INIT_H_DVIN_2B,
      INIT_2C => INIT_H_DVIN_2C,
      INIT_2D => INIT_H_DVIN_2D,
      INIT_2E => INIT_H_DVIN_2E,
      INIT_2F => INIT_H_DVIN_2F,
      INIT_30 => INIT_H_DVIN_30,
      INIT_31 => INIT_H_DVIN_31,
      INIT_32 => INIT_H_DVIN_32,
      INIT_33 => INIT_H_DVIN_33,
      INIT_34 => INIT_H_DVIN_34,
      INIT_35 => INIT_H_DVIN_35,
      INIT_36 => INIT_H_DVIN_36,
      INIT_37 => INIT_H_DVIN_37,
      INIT_38 => INIT_H_DVIN_38,
      INIT_39 => INIT_H_DVIN_39,
      INIT_3A => INIT_H_DVIN_3A,
      INIT_3B => INIT_H_DVIN_3B,
      INIT_3C => INIT_H_DVIN_3C,
      INIT_3D => INIT_H_DVIN_3D,
      INIT_3E => INIT_H_DVIN_3E,
      INIT_3F => INIT_H_DVIN_3F,
      INIT_40 => INIT_H_DVIN_40,
      INIT_41 => INIT_H_DVIN_41,
      INIT_42 => INIT_H_DVIN_42,
      INIT_43 => INIT_H_DVIN_43,
      INIT_44 => INIT_H_DVIN_44,
      INIT_45 => INIT_H_DVIN_45,
      INIT_46 => INIT_H_DVIN_46,
      INIT_47 => INIT_H_DVIN_47,
      INIT_48 => INIT_H_DVIN_48,
      INIT_49 => INIT_H_DVIN_49,
      INIT_4A => INIT_H_DVIN_4A,
      INIT_4B => INIT_H_DVIN_4B,
      INIT_4C => INIT_H_DVIN_4C,
      INIT_4D => INIT_H_DVIN_4D,
      INIT_4E => INIT_H_DVIN_4E,
      INIT_4F => INIT_H_DVIN_4F,
      INIT_50 => INIT_H_DVIN_50,
      INIT_51 => INIT_H_DVIN_51,
      INIT_52 => INIT_H_DVIN_52,
      INIT_53 => INIT_H_DVIN_53,
      INIT_54 => INIT_H_DVIN_54,
      INIT_55 => INIT_H_DVIN_55,
      INIT_56 => INIT_H_DVIN_56,
      INIT_57 => INIT_H_DVIN_57,
      INIT_58 => INIT_H_DVIN_58,
      INIT_59 => INIT_H_DVIN_59,
      INIT_5A => INIT_H_DVIN_5A,
      INIT_5B => INIT_H_DVIN_5B,
      INIT_5C => INIT_H_DVIN_5C,
      INIT_5D => INIT_H_DVIN_5D,
      INIT_5E => INIT_H_DVIN_5E,
      INIT_5F => INIT_H_DVIN_5F,
      INIT_60 => INIT_H_DVIN_60,
      INIT_61 => INIT_H_DVIN_61,
      INIT_62 => INIT_H_DVIN_62,
      INIT_63 => INIT_H_DVIN_63,
      INIT_64 => INIT_H_DVIN_64,
      INIT_65 => INIT_H_DVIN_65,
      INIT_66 => INIT_H_DVIN_66,
      INIT_67 => INIT_H_DVIN_67,
      INIT_68 => INIT_H_DVIN_68,
      INIT_69 => INIT_H_DVIN_69,
      INIT_6A => INIT_H_DVIN_6A,
      INIT_6B => INIT_H_DVIN_6B,
      INIT_6C => INIT_H_DVIN_6C,
      INIT_6D => INIT_H_DVIN_6D,
      INIT_6E => INIT_H_DVIN_6E,
      INIT_6F => INIT_H_DVIN_6F,
      INIT_70 => INIT_H_DVIN_70,
      INIT_71 => INIT_H_DVIN_71,
      INIT_72 => INIT_H_DVIN_72,
      INIT_73 => INIT_H_DVIN_73,
      INIT_74 => INIT_H_DVIN_74,
      INIT_75 => INIT_H_DVIN_75,
      INIT_76 => INIT_H_DVIN_76,
      INIT_77 => INIT_H_DVIN_77,
      INIT_78 => INIT_H_DVIN_78,
      INIT_79 => INIT_H_DVIN_79,
      INIT_7A => INIT_H_DVIN_7A,
      INIT_7B => INIT_H_DVIN_7B,
      INIT_7C => INIT_H_DVIN_7C,
      INIT_7D => INIT_H_DVIN_7D,
      INIT_7E => INIT_H_DVIN_7E,
      INIT_7F => INIT_H_DVIN_7F
   ) port map(
      ADDRARDADDR    => dvin_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => dvin_h_data_out_a(31 downto 0),
      DOPADOP        => dvin_h_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );



   dvin_l_rom: RAMB36E1 generic map (
      READ_WIDTH_A => 9,
      WRITE_WIDTH_A => 9,
      DOA_REG => 0,
      INIT_A => X"000000000",
      RSTREG_PRIORITY_A => "REGCE",
      SRVAL_A => X"000000000",
      WRITE_MODE_A => "WRITE_FIRST",
      READ_WIDTH_B => 9,
      WRITE_WIDTH_B => 9,
      DOB_REG => 0,
      INIT_B => X"000000000",
      RSTREG_PRIORITY_B => "REGCE",
      SRVAL_B => X"000000000",
      WRITE_MODE_B => "WRITE_FIRST",
      INIT_FILE => "NONE",
      SIM_COLLISION_CHECK => "ALL",
      RAM_MODE => "TDP",
      RDADDR_COLLISION_HWCONFIG => "DELAYED_WRITE",
      EN_ECC_READ => FALSE,
      EN_ECC_WRITE => FALSE,
      RAM_EXTENSION_A => "NONE",
      RAM_EXTENSION_B => "NONE",
      SIM_DEVICE => "7SERIES",
      INIT_00 => INIT_L_DVIN_00,
      INIT_01 => INIT_L_DVIN_01,
      INIT_02 => INIT_L_DVIN_02,
      INIT_03 => INIT_L_DVIN_03,
      INIT_04 => INIT_L_DVIN_04,
      INIT_05 => INIT_L_DVIN_05,
      INIT_06 => INIT_L_DVIN_06,
      INIT_07 => INIT_L_DVIN_07,
      INIT_08 => INIT_L_DVIN_08,
      INIT_09 => INIT_L_DVIN_09,
      INIT_0A => INIT_L_DVIN_0A,
      INIT_0B => INIT_L_DVIN_0B,
      INIT_0C => INIT_L_DVIN_0C,
      INIT_0D => INIT_L_DVIN_0D,
      INIT_0E => INIT_L_DVIN_0E,
      INIT_0F => INIT_L_DVIN_0F,
      INIT_10 => INIT_L_DVIN_10,
      INIT_11 => INIT_L_DVIN_11,
      INIT_12 => INIT_L_DVIN_12,
      INIT_13 => INIT_L_DVIN_13,
      INIT_14 => INIT_L_DVIN_14,
      INIT_15 => INIT_L_DVIN_15,
      INIT_16 => INIT_L_DVIN_16,
      INIT_17 => INIT_L_DVIN_17,
      INIT_18 => INIT_L_DVIN_18,
      INIT_19 => INIT_L_DVIN_19,
      INIT_1A => INIT_L_DVIN_1A,
      INIT_1B => INIT_L_DVIN_1B,
      INIT_1C => INIT_L_DVIN_1C,
      INIT_1D => INIT_L_DVIN_1D,
      INIT_1E => INIT_L_DVIN_1E,
      INIT_1F => INIT_L_DVIN_1F,
      INIT_20 => INIT_L_DVIN_20,
      INIT_21 => INIT_L_DVIN_21,
      INIT_22 => INIT_L_DVIN_22,
      INIT_23 => INIT_L_DVIN_23,
      INIT_24 => INIT_L_DVIN_24,
      INIT_25 => INIT_L_DVIN_25,
      INIT_26 => INIT_L_DVIN_26,
      INIT_27 => INIT_L_DVIN_27,
      INIT_28 => INIT_L_DVIN_28,
      INIT_29 => INIT_L_DVIN_29,
      INIT_2A => INIT_L_DVIN_2A,
      INIT_2B => INIT_L_DVIN_2B,
      INIT_2C => INIT_L_DVIN_2C,
      INIT_2D => INIT_L_DVIN_2D,
      INIT_2E => INIT_L_DVIN_2E,
      INIT_2F => INIT_L_DVIN_2F,
      INIT_30 => INIT_L_DVIN_30,
      INIT_31 => INIT_L_DVIN_31,
      INIT_32 => INIT_L_DVIN_32,
      INIT_33 => INIT_L_DVIN_33,
      INIT_34 => INIT_L_DVIN_34,
      INIT_35 => INIT_L_DVIN_35,
      INIT_36 => INIT_L_DVIN_36,
      INIT_37 => INIT_L_DVIN_37,
      INIT_38 => INIT_L_DVIN_38,
      INIT_39 => INIT_L_DVIN_39,
      INIT_3A => INIT_L_DVIN_3A,
      INIT_3B => INIT_L_DVIN_3B,
      INIT_3C => INIT_L_DVIN_3C,
      INIT_3D => INIT_L_DVIN_3D,
      INIT_3E => INIT_L_DVIN_3E,
      INIT_3F => INIT_L_DVIN_3F,
      INIT_40 => INIT_L_DVIN_40,
      INIT_41 => INIT_L_DVIN_41,
      INIT_42 => INIT_L_DVIN_42,
      INIT_43 => INIT_L_DVIN_43,
      INIT_44 => INIT_L_DVIN_44,
      INIT_45 => INIT_L_DVIN_45,
      INIT_46 => INIT_L_DVIN_46,
      INIT_47 => INIT_L_DVIN_47,
      INIT_48 => INIT_L_DVIN_48,
      INIT_49 => INIT_L_DVIN_49,
      INIT_4A => INIT_L_DVIN_4A,
      INIT_4B => INIT_L_DVIN_4B,
      INIT_4C => INIT_L_DVIN_4C,
      INIT_4D => INIT_L_DVIN_4D,
      INIT_4E => INIT_L_DVIN_4E,
      INIT_4F => INIT_L_DVIN_4F,
      INIT_50 => INIT_L_DVIN_50,
      INIT_51 => INIT_L_DVIN_51,
      INIT_52 => INIT_L_DVIN_52,
      INIT_53 => INIT_L_DVIN_53,
      INIT_54 => INIT_L_DVIN_54,
      INIT_55 => INIT_L_DVIN_55,
      INIT_56 => INIT_L_DVIN_56,
      INIT_57 => INIT_L_DVIN_57,
      INIT_58 => INIT_L_DVIN_58,
      INIT_59 => INIT_L_DVIN_59,
      INIT_5A => INIT_L_DVIN_5A,
      INIT_5B => INIT_L_DVIN_5B,
      INIT_5C => INIT_L_DVIN_5C,
      INIT_5D => INIT_L_DVIN_5D,
      INIT_5E => INIT_L_DVIN_5E,
      INIT_5F => INIT_L_DVIN_5F,
      INIT_60 => INIT_L_DVIN_60,
      INIT_61 => INIT_L_DVIN_61,
      INIT_62 => INIT_L_DVIN_62,
      INIT_63 => INIT_L_DVIN_63,
      INIT_64 => INIT_L_DVIN_64,
      INIT_65 => INIT_L_DVIN_65,
      INIT_66 => INIT_L_DVIN_66,
      INIT_67 => INIT_L_DVIN_67,
      INIT_68 => INIT_L_DVIN_68,
      INIT_69 => INIT_L_DVIN_69,
      INIT_6A => INIT_L_DVIN_6A,
      INIT_6B => INIT_L_DVIN_6B,
      INIT_6C => INIT_L_DVIN_6C,
      INIT_6D => INIT_L_DVIN_6D,
      INIT_6E => INIT_L_DVIN_6E,
      INIT_6F => INIT_L_DVIN_6F,
      INIT_70 => INIT_L_DVIN_70,
      INIT_71 => INIT_L_DVIN_71,
      INIT_72 => INIT_L_DVIN_72,
      INIT_73 => INIT_L_DVIN_73,
      INIT_74 => INIT_L_DVIN_74,
      INIT_75 => INIT_L_DVIN_75,
      INIT_76 => INIT_L_DVIN_76,
      INIT_77 => INIT_L_DVIN_77,
      INIT_78 => INIT_L_DVIN_78,
      INIT_79 => INIT_L_DVIN_79,
      INIT_7A => INIT_L_DVIN_7A,
      INIT_7B => INIT_L_DVIN_7B,
      INIT_7C => INIT_L_DVIN_7C,
      INIT_7D => INIT_L_DVIN_7D,
      INIT_7E => INIT_L_DVIN_7E,
      INIT_7F => INIT_L_DVIN_7F
   ) port map(
      ADDRARDADDR    => dvin_address_a,
      ENARDEN        => '1',
      CLKARDCLK      => sysClk,
      DOADO          => dvin_l_data_out_a(31 downto 0),
      DOPADOP        => dvin_l_data_out_a(35 downto 32),
      DIADI          => x"00000000",
      DIPADIP        => x"0",
      WEA            => "0000",
      REGCEAREGCE    => '0',
      RSTRAMARSTRAM  => '0',
      RSTREGARSTREG  => '0',
      ADDRBWRADDR    => x"0000",
      ENBWREN        => '0',
      CLKBWRCLK      => sysClk,
      DOBDO          => open,
      DOPBDOP        => open,
      DIBDI          => x"00000000",
      DIPBDIP        => x"0",
      WEBWE          => x"00",
      REGCEB         => '0',
      RSTRAMB        => '0',
      RSTREGB        => '0',
      CASCADEINA     => '0',
      CASCADEINB     => '0',
      INJECTDBITERR  => '0',
      INJECTSBITERR  => '0'
   );

   dvin_address_a <= '1' & adcData(8)(23 downto 12) & "111";
   outEnvData(8) <= x"0000" & dvin_h_data_out_a(7 downto 0) & dvin_l_data_out_a(7 downto 0);

end RTL;

